(**
  This file defines the meta-level functions to express the module system of
  (Core) Erlang.
*)

From CoreErlang.BigStep Require Export Auxiliaries.

Import ListNotations.

(* Module Helpers with records *)
Fixpoint get_module (name' : string) (ml : list ErlModule) : option ErlModule := 
    match ml with
    | m :: ms => if (eqb  (name m)  name')  then Some m else get_module name' ms
    | [] => None
end
.

(* Checks if a function is in the list of function identifiers*)
Fixpoint check_in_functions (name : string) (arity : nat) (fl: list FunctionIdentifier) : bool :=
    match fl with
    | f :: fs => if 
                    andb 
                      (eqb (fst f) name) 
                      (Nat.eqb (snd f) arity)
                    then
                      true
                    else
                      check_in_functions name arity fs 
    | [] => false
end.

(* Returns a function from a list of top-level function by name *)
Fixpoint get_function (name : string) (arity : nat) (fl: list TopLevelFunction) : option TopLevelFunction:=
    match fl with
    | f :: fs => if andb 
                      (eqb (fst (identifier f)) (name)) 
                      (Nat.eqb (snd (identifier f)) (arity))
                  then
                    Some f 
                  else
                    get_function name arity fs
    | [] => None
end.

Definition get_modfunc (mname : string) (fname : string) (arity : nat) (ml : list ErlModule) : option TopLevelFunction  :=
    match get_module mname ml with
    | Some m => 
        if check_in_functions fname arity (funcIds m) then
                get_function fname arity (funcs m)
            else
                None
    | None => None
end.

Definition get_own_modfunc (mname : string) (fname : string) (arity : nat) (ml : list ErlModule) : option TopLevelFunction  :=
    match get_module mname ml with
    | Some m => get_function fname arity (funcs m)
    | None => None
end.



(* Standard library *)
Definition stdlib : list ErlModule :=
  [
    (* Lists module*)
    {| 
      name := "lists"%string;
      funcIds := [
          ("all"%string, 2);("any"%string, 2);
          ("append"%string, 1);
          ("append"%string, 2);
          ("concat"%string, 1);
          ("delete"%string, 2);
          ("droplast"%string, 1);
          ("dropwhile"%string, 2);
          ("duplicate"%string, 2);
          ("enumerate"%string, 1);
          ("enumerate"%string, 2);
          ("filter"%string, 2);
          ("filtermap"%string, 2);
          ("flatlength"%string, 1);
          ("flatmap"%string, 2);
          ("flatten"%string, 1);
          ("flatten"%string, 2);
          ("foldl"%string, 3);
          ("foldr"%string, 3);
          ("foreach"%string, 2);
          ("join"%string, 2);
          ("keydelete"%string, 3);
          ("keyfind"%string, 3);
          ("keymap"%string, 3);
          ("keymember"%string, 3);
          ("keymerge"%string, 3);
          ("keyreplace"%string, 4);
          ("keysearch"%string, 3);
          ("keysort"%string, 2);
          ("keystore"%string, 4);
          ("keytake"%string, 3);
          ("last"%string, 1);
          ("map"%string, 2);
          ("mapfoldl"%string, 3);
          ("mapfoldr"%string, 3);
          ("max"%string, 1);
          ("member"%string, 2);
          ("merge"%string, 1);
          ("merge"%string, 2);
          ("merge"%string, 3);
          ("merge3"%string, 3);
          ("min"%string, 1);
          ("module_info"%string, 0);
          ("module_info"%string, 1);
          ("nth"%string, 2);
          ("nthtail"%string, 2);
          ("partition"%string, 2);
          ("prefix"%string, 2);
          ("reverse"%string, 1);
          ("reverse"%string, 2);
          ("rkeymerge"%string, 3);
          ("rmerge"%string, 2);
          ("rmerge"%string, 3);
          ("rmerge3"%string, 3);
          ("rukeymerge"%string, 3);
          ("rumerge"%string, 2);
          ("rumerge"%string, 3);
          ("rumerge3"%string, 3);
          ("search"%string, 2);
          ("seq"%string, 2);
          ("seq"%string, 3);
          ("sort"%string, 1);
          ("sort"%string, 2);
          ("split"%string, 2);
          ("splitwith"%string, 2);
          ("sublist"%string, 2);
          ("sublist"%string, 3);
          ("subtract"%string, 2);
          ("suffix"%string, 2);
          ("sum"%string, 1);
          ("takewhile"%string, 2);
          ("ukeymerge"%string, 3);
          ("ukeysort"%string, 2);
          ("umerge"%string, 1);
          ("umerge"%string, 2);
          ("umerge"%string, 3);
          ("umerge3"%string, 3);
          ("uniq"%string, 1);
          ("uniq"%string, 2);
          ("unzip"%string, 1);
          ("unzip3"%string, 1);
          ("usort"%string, 1);
          ("usort"%string, 2);
          ("zf"%string, 2);
          ("zip"%string, 2);
          ("zip3"%string, 3);
          ("zipwith"%string, 3);
          ("zipwith3"%string, 4)];
      attrs := []; 
      funcs := [
          {| identifier := ("keyfind"%string, 3) ; varl := ["_0"%string;"_1"%string;"_2"%string]; body := (ECase (EApp (EFunId ("keysearch"%string, 3)) [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string)]) [([(PTuple [(PVar "_7"%string);(PVar "Tuple"%string)])], (ELit (Atom "true"%string)), (EVar "Tuple"%string));([(PVar "X"%string)], (ELit (Atom "true"%string)), (EVar "X"%string))]) |};
          {| identifier := ("keymember"%string, 3) ; varl := ["_0"%string;"_1"%string;"_2"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string)]) [([(PVar "K"%string);(PVar "N"%string);(PVar "L"%string)], (ELet ["_3"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_integer"%string)) [(EVar "N"%string)]) (ELet ["_4"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom ">"%string)) [(EVar "N"%string);(ELit (Integer (0)))]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "and"%string)) [(EVar "_3"%string);(EVar "_4"%string)]))), (EApp (EFunId ("keymember3"%string, 3)) [(EVar "K"%string);(EVar "N"%string);(EVar "L"%string)]));([(PVar "_7"%string);(PVar "_6"%string);(PVar "_5"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_7"%string);(EVar "_6"%string);(EVar "_5"%string)])]))]) |};
          {| identifier := ("keymember3"%string, 3) ; varl := ["_0"%string;"_1"%string;"_2"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string)]) [([(PVar "Key"%string);(PVar "N"%string);(PCons (PVar "T"%string) (PVar "Ts"%string))], (ETry (ELet ["_3"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "N"%string);(EVar "T"%string)]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "_3"%string);(EVar "Key"%string)])) ["Try"%string] (EVar "Try"%string) ["T"%string;"R"%string] (ELit (Atom "false"%string))), (ELit (Atom "true"%string)));([(PVar "Key"%string);(PVar "N"%string);(PCons (PVar "T"%string) (PVar "Ts"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("keymember3"%string, 3)) [(EVar "Key"%string);(EVar "N"%string);(EVar "Ts"%string)]));([(PVar "Key"%string);(PVar "N"%string);PNil], (ELit (Atom "true"%string)), (ELit (Atom "false"%string)));([(PVar "_6"%string);(PVar "_5"%string);(PVar "_4"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_6"%string);(EVar "_5"%string);(EVar "_4"%string)])]))]) |};
          {| identifier := ("keysearch"%string, 3) ; varl := ["_0"%string;"_1"%string;"_2"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string)]) [([(PVar "K"%string);(PVar "N"%string);(PVar "L"%string)], (ELet ["_3"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_integer"%string)) [(EVar "N"%string)]) (ELet ["_4"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom ">"%string)) [(EVar "N"%string);(ELit (Integer (0)))]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "and"%string)) [(EVar "_3"%string);(EVar "_4"%string)]))), (EApp (EFunId ("keysearch3"%string, 3)) [(EVar "K"%string);(EVar "N"%string);(EVar "L"%string)]));([(PVar "_7"%string);(PVar "_6"%string);(PVar "_5"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_7"%string);(EVar "_6"%string);(EVar "_5"%string)])]))]) |};
          {| identifier := ("keysearch3"%string, 3) ; varl := ["_0"%string;"_1"%string;"_2"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string)]) [([(PVar "Key"%string);(PVar "N"%string);(PCons (PVar "H"%string) (PVar "T"%string))], (ETry (ELet ["_3"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "N"%string);(EVar "H"%string)]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "_3"%string);(EVar "Key"%string)])) ["Try"%string] (EVar "Try"%string) ["T"%string;"R"%string] (ELit (Atom "false"%string))), (ETuple [(ELit (Atom "value"%string));(EVar "H"%string)]));([(PVar "Key"%string);(PVar "N"%string);(PCons (PVar "H"%string) (PVar "T"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("keysearch3"%string, 3)) [(EVar "Key"%string);(EVar "N"%string);(EVar "T"%string)]));([(PVar "Key"%string);(PVar "N"%string);PNil], (ELit (Atom "true"%string)), (ELit (Atom "false"%string)));([(PVar "_6"%string);(PVar "_5"%string);(PVar "_4"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_6"%string);(EVar "_5"%string);(EVar "_4"%string)])]))]) |};
          {| identifier := ("member"%string, 2) ; varl := ["_0"%string;"_1"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string)]) [([(PVar "X"%string);(PCons (PVar "_4"%string) (PVar "_5"%string))], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=:="%string)) [(EVar "_4"%string);(EVar "X"%string)]), (ELit (Atom "true"%string)));([(PVar "X"%string);(PCons (PVar "_6"%string) (PVar "Y"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("member"%string, 2)) [(EVar "X"%string);(EVar "Y"%string)]));([(PVar "X"%string);PNil], (ELit (Atom "true"%string)), (ELit (Atom "false"%string)));([(PVar "_3"%string);(PVar "_2"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_3"%string);(EVar "_2"%string)])]))]) |};
          {| identifier := ("reverse"%string, 2) ; varl := ["_0"%string;"_1"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string)]) [([(PCons (PVar "H"%string) (PVar "T"%string));(PVar "Y"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("reverse"%string, 2)) [(EVar "T"%string);(ECons (EVar "H"%string) (EVar "Y"%string))]));([PNil;(PVar "X"%string)], (ELit (Atom "true"%string)), (EVar "X"%string));([(PVar "_3"%string);(PVar "_2"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_3"%string);(EVar "_2"%string)])]))]) |};
          {| identifier := ("append"%string, 2) ; varl := ["_0"%string;"_1"%string]; body := (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "++"%string)) [(EVar "_0"%string);(EVar "_1"%string)]) |};
          {| identifier := ("append"%string, 1) ; varl := ["_0"%string]; body := (ECase (EVar "_0"%string) [([(PCons (PVar "E"%string) PNil)], (ELit (Atom "true"%string)), (EVar "E"%string));([(PCons (PVar "H"%string) (PVar "T"%string))], (ELit (Atom "true"%string)), (ELet ["_1"%string] (EApp (EFunId ("append"%string, 1)) [(EVar "T"%string)]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "++"%string)) [(EVar "H"%string);(EVar "_1"%string)])));([PNil], (ELit (Atom "true"%string)), ENil);([(PVar "_2"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_2"%string)])]))]) |};
          {| identifier := ("subtract"%string, 2) ; varl := ["_0"%string;"_1"%string]; body := (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "--"%string)) [(EVar "_0"%string);(EVar "_1"%string)]) |};
          {| identifier := ("reverse"%string, 1) ; varl := ["_0"%string]; body := (ECase (EVar "_0"%string) [([(PTuple [(PLit (Atom "c_alias"%string));PNil;(PVar "L"%string);PNil])], (ELit (Atom "true"%string)), (EVar "L"%string));([(PTuple [(PLit (Atom "c_alias"%string));PNil;(PVar "L"%string);(PCons (PVar "_2"%string) PNil)])], (ELit (Atom "true"%string)), (EVar "L"%string));([(PCons (PVar "A"%string) (PCons (PVar "B"%string) PNil))], (ELit (Atom "true"%string)), (ECons (EVar "B"%string) (ECons (EVar "A"%string) ENil)));([(PCons (PVar "A"%string) (PCons (PVar "B"%string) (PVar "L"%string)))], (ELit (Atom "true"%string)), (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "L"%string);(ECons (EVar "B"%string) (ECons (EVar "A"%string) ENil))]));([(PVar "_1"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_1"%string)])]))]) |};
          {| identifier := ("nth"%string, 2) ; varl := ["_0"%string;"_1"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string)]) [([(PLit (Integer (1)));(PCons (PVar "H"%string) (PVar "_5"%string))], (ELit (Atom "true"%string)), (EVar "H"%string));([(PVar "N"%string);(PCons (PVar "_6"%string) (PVar "T"%string))], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom ">"%string)) [(EVar "N"%string);(ELit (Integer (1)))]), (ELet ["_2"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "-"%string)) [(EVar "N"%string);(ELit (Integer (1)))]) (EApp (EFunId ("nth"%string, 2)) [(EVar "_2"%string);(EVar "T"%string)])));([(PVar "_4"%string);(PVar "_3"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_4"%string);(EVar "_3"%string)])]))]) |};
          {| identifier := ("nthtail"%string, 2) ; varl := ["_0"%string;"_1"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string)]) [([(PLit (Integer (1)));(PCons (PVar "_5"%string) (PVar "T"%string))], (ELit (Atom "true"%string)), (EVar "T"%string));([(PVar "N"%string);(PCons (PVar "_6"%string) (PVar "T"%string))], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom ">"%string)) [(EVar "N"%string);(ELit (Integer (1)))]), (ELet ["_2"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "-"%string)) [(EVar "N"%string);(ELit (Integer (1)))]) (EApp (EFunId ("nthtail"%string, 2)) [(EVar "_2"%string);(EVar "T"%string)])));([(PLit (Integer (0)));(PVar "L"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_list"%string)) [(EVar "L"%string)]), (EVar "L"%string));([(PVar "_4"%string);(PVar "_3"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_4"%string);(EVar "_3"%string)])]))]) |};
          {| identifier := ("prefix"%string, 2) ; varl := ["_0"%string;"_1"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string)]) [([(PCons (PVar "X"%string) (PVar "PreTail"%string));(PCons (PVar "_4"%string) (PVar "Tail"%string))], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=:="%string)) [(EVar "_4"%string);(EVar "X"%string)]), (EApp (EFunId ("prefix"%string, 2)) [(EVar "PreTail"%string);(EVar "Tail"%string)]));([PNil;(PVar "List"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_list"%string)) [(EVar "List"%string)]), (ELit (Atom "true"%string)));([(PCons (PVar "_5"%string) (PVar "_6"%string));(PVar "List"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_list"%string)) [(EVar "List"%string)]), (ELit (Atom "false"%string)));([(PVar "_3"%string);(PVar "_2"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_3"%string);(EVar "_2"%string)])]))]) |};
          {| identifier := ("suffix"%string, 2) ; varl := ["_0"%string;"_1"%string]; body := (ELet ["_3"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "length"%string)) [(EVar "_1"%string)]) (ELet ["_2"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "length"%string)) [(EVar "_0"%string)]) (ELet ["Delta"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "-"%string)) [(EVar "_3"%string);(EVar "_2"%string)]) (ECase (ECall (ELit (Atom "erlang"%string)) (ELit (Atom ">="%string)) [(EVar "Delta"%string);(ELit (Integer (0)))]) [([(PLit (Atom "true"%string))], (ELit (Atom "true"%string)), (ELet ["_6"%string] (EApp (EFunId ("nthtail"%string, 2)) [(EVar "Delta"%string);(EVar "_1"%string)]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=:="%string)) [(EVar "_6"%string);(EVar "_0"%string)])));([(PLit (Atom "false"%string))], (ELit (Atom "true"%string)), (ELit (Atom "false"%string)))])))) |};
          {| identifier := ("droplast"%string, 1) ; varl := ["_0"%string]; body := (ECase (EVar "_0"%string) [([(PCons (PVar "_T"%string) PNil)], (ELit (Atom "true"%string)), ENil);([(PCons (PVar "H"%string) (PVar "T"%string))], (ELit (Atom "true"%string)), (ELet ["_1"%string] (EApp (EFunId ("droplast"%string, 1)) [(EVar "T"%string)]) (ECons (EVar "H"%string) (EVar "_1"%string))));([(PVar "_2"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_2"%string)])]))]) |};
          {| identifier := ("last"%string, 1) ; varl := ["_0"%string]; body := (ECase (EVar "_0"%string) [([(PCons (PVar "E"%string) (PVar "Es"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("last"%string, 2)) [(EVar "E"%string);(EVar "Es"%string)]));([(PVar "_1"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_1"%string)])]))]) |};
          {| identifier := ("last"%string, 2) ; varl := ["_0"%string;"_1"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string)]) [([(PVar "_4"%string);(PCons (PVar "E"%string) (PVar "Es"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("last"%string, 2)) [(EVar "E"%string);(EVar "Es"%string)]));([(PVar "E"%string);PNil], (ELit (Atom "true"%string)), (EVar "E"%string));([(PVar "_3"%string);(PVar "_2"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_3"%string);(EVar "_2"%string)])]))]) |};
          {| identifier := ("seq"%string, 2) ; varl := ["_0"%string;"_1"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string)]) [([(PVar "First"%string);(PVar "Last"%string)], (ETry (ELet ["_2"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_integer"%string)) [(EVar "First"%string)]) (ELet ["_3"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_integer"%string)) [(EVar "Last"%string)]) (ELet ["_4"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "-"%string)) [(EVar "First"%string);(ELit (Integer (1)))]) (ELet ["_5"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "_4"%string);(EVar "Last"%string)]) (ELet ["_6"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "and"%string)) [(EVar "_3"%string);(EVar "_5"%string)]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "and"%string)) [(EVar "_2"%string);(EVar "_6"%string)])))))) ["Try"%string] (EVar "Try"%string) ["T"%string;"R"%string] (ELit (Atom "false"%string))), (ELet ["_7"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "-"%string)) [(EVar "Last"%string);(EVar "First"%string)]) (ELet ["_8"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "+"%string)) [(EVar "_7"%string);(ELit (Integer (1)))]) (EApp (EFunId ("seq_loop"%string, 3)) [(EVar "_8"%string);(EVar "Last"%string);ENil]))));([(PVar "_10"%string);(PVar "_9"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_10"%string);(EVar "_9"%string)])]))]) |};
          {| identifier := ("seq_loop"%string, 3) ; varl := ["_0"%string;"_1"%string;"_2"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string)]) [([(PVar "N"%string);(PVar "X"%string);(PVar "L"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom ">="%string)) [(EVar "N"%string);(ELit (Integer (4)))]), (ELet ["_7"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "-"%string)) [(EVar "N"%string);(ELit (Integer (4)))]) (ELet ["_6"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "-"%string)) [(EVar "X"%string);(ELit (Integer (4)))]) (ELet ["_3"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "-"%string)) [(EVar "X"%string);(ELit (Integer (3)))]) (ELet ["_4"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "-"%string)) [(EVar "X"%string);(ELit (Integer (2)))]) (ELet ["_5"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "-"%string)) [(EVar "X"%string);(ELit (Integer (1)))]) (EApp (EFunId ("seq_loop"%string, 3)) [(EVar "_7"%string);(EVar "_6"%string);(ECons (EVar "_3"%string) (ECons (EVar "_4"%string) (ECons (EVar "_5"%string) (ECons (EVar "X"%string) (EVar "L"%string)))))])))))));([(PVar "N"%string);(PVar "X"%string);(PVar "L"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom ">="%string)) [(EVar "N"%string);(ELit (Integer (2)))]), (ELet ["_10"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "-"%string)) [(EVar "N"%string);(ELit (Integer (2)))]) (ELet ["_9"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "-"%string)) [(EVar "X"%string);(ELit (Integer (2)))]) (ELet ["_8"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "-"%string)) [(EVar "X"%string);(ELit (Integer (1)))]) (EApp (EFunId ("seq_loop"%string, 3)) [(EVar "_10"%string);(EVar "_9"%string);(ECons (EVar "_8"%string) (ECons (EVar "X"%string) (EVar "L"%string)))])))));([(PLit (Integer (1)));(PVar "X"%string);(PVar "L"%string)], (ELit (Atom "true"%string)), (ECons (EVar "X"%string) (EVar "L"%string)));([(PLit (Integer (0)));(PVar "_14"%string);(PVar "L"%string)], (ELit (Atom "true"%string)), (EVar "L"%string));([(PVar "_13"%string);(PVar "_12"%string);(PVar "_11"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_13"%string);(EVar "_12"%string);(EVar "_11"%string)])]))]) |};
          {| identifier := ("seq"%string, 3) ; varl := ["_0"%string;"_1"%string;"_2"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string)]) [([(PVar "First"%string);(PVar "Last"%string);(PVar "Inc"%string)], (ETry (ELet ["_3"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_integer"%string)) [(EVar "First"%string)]) (ELet ["_4"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_integer"%string)) [(EVar "Last"%string)]) (ELet ["_5"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_integer"%string)) [(EVar "Inc"%string)]) (ELet ["_10"%string] (ECase (ECall (ELit (Atom "erlang"%string)) (ELit (Atom ">"%string)) [(EVar "Inc"%string);(ELit (Integer (0)))]) [([(PLit (Atom "true"%string))], (ELit (Atom "true"%string)), (ELet ["_8"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "-"%string)) [(EVar "First"%string);(EVar "Inc"%string)]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "_8"%string);(EVar "Last"%string)])));([(PLit (Atom "false"%string))], (ELit (Atom "true"%string)), (ELit (Atom "false"%string)));([(PVar "_7"%string)], (ELit (Atom "true"%string)), (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "error"%string)) [(ETuple [(ELit (Atom "badarg"%string));(EVar "_7"%string)])]))]) (ELet ["_15"%string] (ECase (EVar "_10"%string) [([(PLit (Atom "true"%string))], (ELit (Atom "true"%string)), (ELit (Atom "true"%string)));([(PLit (Atom "false"%string))], (ELit (Atom "true"%string)), (ECase (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "<"%string)) [(EVar "Inc"%string);(ELit (Integer (0)))]) [([(PLit (Atom "true"%string))], (ELit (Atom "true"%string)), (ELet ["_12"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "-"%string)) [(EVar "First"%string);(EVar "Inc"%string)]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom ">="%string)) [(EVar "_12"%string);(EVar "Last"%string)])));([(PLit (Atom "false"%string))], (ELit (Atom "true"%string)), (ELit (Atom "false"%string)));([(PVar "_11"%string)], (ELit (Atom "true"%string)), (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "error"%string)) [(ETuple [(ELit (Atom "badarg"%string));(EVar "_11"%string)])]))]));([(PVar "_6"%string)], (ELit (Atom "true"%string)), (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "error"%string)) [(ETuple [(ELit (Atom "badarg"%string));(EVar "_6"%string)])]))]) (ELet ["_16"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=:="%string)) [(EVar "_15"%string);(ELit (Atom "true"%string))]) (ELet ["_17"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "and"%string)) [(EVar "_5"%string);(EVar "_16"%string)]) (ELet ["_18"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "and"%string)) [(EVar "_4"%string);(EVar "_17"%string)]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "and"%string)) [(EVar "_3"%string);(EVar "_18"%string)]))))))))) ["Try"%string] (EVar "Try"%string) ["T"%string;"R"%string] (ELit (Atom "false"%string))), (ELet ["_19"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "-"%string)) [(EVar "Last"%string);(EVar "First"%string)]) (ELet ["_20"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "+"%string)) [(EVar "_19"%string);(EVar "Inc"%string)]) (ELet ["N"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "div"%string)) [(EVar "_20"%string);(EVar "Inc"%string)]) (ELet ["_22"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "-"%string)) [(EVar "N"%string);(ELit (Integer (1)))]) (ELet ["_23"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "*"%string)) [(EVar "Inc"%string);(EVar "_22"%string)]) (ELet ["_24"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "+"%string)) [(EVar "_23"%string);(EVar "First"%string)]) (EApp (EFunId ("seq_loop"%string, 4)) [(EVar "N"%string);(EVar "_24"%string);(EVar "Inc"%string);ENil]))))))));([(PVar "Same"%string);(PVar "_28"%string);(PLit (Integer (0)))], (ELet ["_29"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=:="%string)) [(EVar "_28"%string);(EVar "Same"%string)]) (ELet ["_30"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_integer"%string)) [(EVar "Same"%string)]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "and"%string)) [(EVar "_29"%string);(EVar "_30"%string)]))), (ECons (EVar "Same"%string) ENil));([(PVar "First"%string);(PVar "Last"%string);(PVar "Inc"%string)], (ELit (Atom "true"%string)), (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "error"%string)) [(ELit (Atom "badarg"%string));(ECons (EVar "First"%string) (ECons (EVar "Last"%string) (ECons (EVar "Inc"%string) ENil)));(ECons (ETuple [(ELit (Atom "error_info"%string));(EMap [((ELit (Atom "module"%string)),(ELit (Atom "erl_stdlib_errors"%string)))])]) ENil)]))]) |};
          {| identifier := ("seq_loop"%string, 4) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string)]) [([(PVar "N"%string);(PVar "X"%string);(PVar "D"%string);(PVar "L"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom ">="%string)) [(EVar "N"%string);(ELit (Integer (4)))]), (ELet ["Y"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "-"%string)) [(EVar "X"%string);(EVar "D"%string)]) (ELet ["Z"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "-"%string)) [(EVar "Y"%string);(EVar "D"%string)]) (ELet ["W"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "-"%string)) [(EVar "Z"%string);(EVar "D"%string)]) (ELet ["_8"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "-"%string)) [(EVar "N"%string);(ELit (Integer (4)))]) (ELet ["_7"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "-"%string)) [(EVar "W"%string);(EVar "D"%string)]) (EApp (EFunId ("seq_loop"%string, 4)) [(EVar "_8"%string);(EVar "_7"%string);(EVar "D"%string);(ECons (EVar "W"%string) (ECons (EVar "Z"%string) (ECons (EVar "Y"%string) (ECons (EVar "X"%string) (EVar "L"%string)))))])))))));([(PVar "N"%string);(PVar "X"%string);(PVar "D"%string);(PVar "L"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom ">="%string)) [(EVar "N"%string);(ELit (Integer (2)))]), (ELet ["Y"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "-"%string)) [(EVar "X"%string);(EVar "D"%string)]) (ELet ["_11"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "-"%string)) [(EVar "N"%string);(ELit (Integer (2)))]) (ELet ["_10"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "-"%string)) [(EVar "Y"%string);(EVar "D"%string)]) (EApp (EFunId ("seq_loop"%string, 4)) [(EVar "_11"%string);(EVar "_10"%string);(EVar "D"%string);(ECons (EVar "Y"%string) (ECons (EVar "X"%string) (EVar "L"%string)))])))));([(PLit (Integer (1)));(PVar "X"%string);(PVar "_16"%string);(PVar "L"%string)], (ELit (Atom "true"%string)), (ECons (EVar "X"%string) (EVar "L"%string)));([(PLit (Integer (0)));(PVar "_17"%string);(PVar "_18"%string);(PVar "L"%string)], (ELit (Atom "true"%string)), (EVar "L"%string));([(PVar "_15"%string);(PVar "_14"%string);(PVar "_13"%string);(PVar "_12"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_15"%string);(EVar "_14"%string);(EVar "_13"%string);(EVar "_12"%string)])]))]) |};
          {| identifier := ("sum"%string, 1) ; varl := ["_0"%string]; body := (EApp (EFunId ("sum"%string, 2)) [(EVar "_0"%string);(ELit (Integer (0)))]) |};
          {| identifier := ("sum"%string, 2) ; varl := ["_0"%string;"_1"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string)]) [([(PCons (PVar "H"%string) (PVar "T"%string));(PVar "Sum"%string)], (ELit (Atom "true"%string)), (ELet ["_2"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "+"%string)) [(EVar "Sum"%string);(EVar "H"%string)]) (EApp (EFunId ("sum"%string, 2)) [(EVar "T"%string);(EVar "_2"%string)])));([PNil;(PVar "Sum"%string)], (ELit (Atom "true"%string)), (EVar "Sum"%string));([(PVar "_4"%string);(PVar "_3"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_4"%string);(EVar "_3"%string)])]))]) |};
          {| identifier := ("duplicate"%string, 2) ; varl := ["_0"%string;"_1"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string)]) [([(PVar "N"%string);(PVar "X"%string)], (ELet ["_2"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_integer"%string)) [(EVar "N"%string)]) (ELet ["_3"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom ">="%string)) [(EVar "N"%string);(ELit (Integer (0)))]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "and"%string)) [(EVar "_2"%string);(EVar "_3"%string)]))), (EApp (EFunId ("duplicate"%string, 3)) [(EVar "N"%string);(EVar "X"%string);ENil]));([(PVar "_5"%string);(PVar "_4"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_5"%string);(EVar "_4"%string)])]))]) |};
          {| identifier := ("duplicate"%string, 3) ; varl := ["_0"%string;"_1"%string;"_2"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string)]) [([(PLit (Integer (0)));(PVar "_7"%string);(PVar "L"%string)], (ELit (Atom "true"%string)), (EVar "L"%string));([(PVar "N"%string);(PVar "X"%string);(PVar "L"%string)], (ELit (Atom "true"%string)), (ELet ["_3"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "-"%string)) [(EVar "N"%string);(ELit (Integer (1)))]) (EApp (EFunId ("duplicate"%string, 3)) [(EVar "_3"%string);(EVar "X"%string);(ECons (EVar "X"%string) (EVar "L"%string))])))]) |};
          {| identifier := ("min"%string, 1) ; varl := ["_0"%string]; body := (ECase (EVar "_0"%string) [([(PCons (PVar "H"%string) (PVar "T"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("min"%string, 2)) [(EVar "T"%string);(EVar "H"%string)]));([(PVar "_1"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_1"%string)])]))]) |};
          {| identifier := ("min"%string, 2) ; varl := ["_0"%string;"_1"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string)]) [([(PCons (PVar "H"%string) (PVar "T"%string));(PVar "Min"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "<"%string)) [(EVar "H"%string);(EVar "Min"%string)]), (EApp (EFunId ("min"%string, 2)) [(EVar "T"%string);(EVar "H"%string)]));([(PCons (PVar "_4"%string) (PVar "T"%string));(PVar "Min"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("min"%string, 2)) [(EVar "T"%string);(EVar "Min"%string)]));([PNil;(PVar "Min"%string)], (ELit (Atom "true"%string)), (EVar "Min"%string));([(PVar "_3"%string);(PVar "_2"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_3"%string);(EVar "_2"%string)])]))]) |};
          {| identifier := ("max"%string, 1) ; varl := ["_0"%string]; body := (ECase (EVar "_0"%string) [([(PCons (PVar "H"%string) (PVar "T"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("max"%string, 2)) [(EVar "T"%string);(EVar "H"%string)]));([(PVar "_1"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_1"%string)])]))]) |};
          {| identifier := ("max"%string, 2) ; varl := ["_0"%string;"_1"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string)]) [([(PCons (PVar "H"%string) (PVar "T"%string));(PVar "Max"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom ">"%string)) [(EVar "H"%string);(EVar "Max"%string)]), (EApp (EFunId ("max"%string, 2)) [(EVar "T"%string);(EVar "H"%string)]));([(PCons (PVar "_4"%string) (PVar "T"%string));(PVar "Max"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("max"%string, 2)) [(EVar "T"%string);(EVar "Max"%string)]));([PNil;(PVar "Max"%string)], (ELit (Atom "true"%string)), (EVar "Max"%string));([(PVar "_3"%string);(PVar "_2"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_3"%string);(EVar "_2"%string)])]))]) |};
          {| identifier := ("sublist"%string, 3) ; varl := ["_0"%string;"_1"%string;"_2"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string)]) [([(PVar "List"%string);(PLit (Integer (1)));(PVar "L"%string)], (ETry (ELet ["_3"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_list"%string)) [(EVar "List"%string)]) (ELet ["_4"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_integer"%string)) [(EVar "L"%string)]) (ELet ["_5"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom ">="%string)) [(EVar "L"%string);(ELit (Integer (0)))]) (ELet ["_6"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "and"%string)) [(EVar "_4"%string);(EVar "_5"%string)]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "and"%string)) [(EVar "_3"%string);(EVar "_6"%string)]))))) ["Try"%string] (EVar "Try"%string) ["T"%string;"R"%string] (ELit (Atom "false"%string))), (EApp (EFunId ("sublist"%string, 2)) [(EVar "List"%string);(EVar "L"%string)]));([PNil;(PVar "S"%string);(PVar "_L"%string)], (ELet ["_7"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_integer"%string)) [(EVar "S"%string)]) (ELet ["_8"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom ">="%string)) [(EVar "S"%string);(ELit (Integer (2)))]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "and"%string)) [(EVar "_7"%string);(EVar "_8"%string)]))), ENil);([(PCons (PVar "_H"%string) (PVar "T"%string));(PVar "S"%string);(PVar "L"%string)], (ELet ["_9"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_integer"%string)) [(EVar "S"%string)]) (ELet ["_10"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom ">="%string)) [(EVar "S"%string);(ELit (Integer (2)))]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "and"%string)) [(EVar "_9"%string);(EVar "_10"%string)]))), (ELet ["_11"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "-"%string)) [(EVar "S"%string);(ELit (Integer (1)))]) (EApp (EFunId ("sublist"%string, 3)) [(EVar "T"%string);(EVar "_11"%string);(EVar "L"%string)])));([(PVar "_14"%string);(PVar "_13"%string);(PVar "_12"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_14"%string);(EVar "_13"%string);(EVar "_12"%string)])]))]) |};
          {| identifier := ("sublist"%string, 2) ; varl := ["_0"%string;"_1"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string)]) [([(PVar "List"%string);(PVar "L"%string)], (ELet ["_2"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_integer"%string)) [(EVar "L"%string)]) (ELet ["_3"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_list"%string)) [(EVar "List"%string)]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "and"%string)) [(EVar "_2"%string);(EVar "_3"%string)]))), (EApp (EFunId ("sublist_2"%string, 2)) [(EVar "List"%string);(EVar "L"%string)]));([(PVar "_5"%string);(PVar "_4"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_5"%string);(EVar "_4"%string)])]))]) |};
          {| identifier := ("sublist_2"%string, 2) ; varl := ["_0"%string;"_1"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string)]) [([(PCons (PVar "H"%string) (PVar "T"%string));(PVar "L"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom ">"%string)) [(EVar "L"%string);(ELit (Integer (0)))]), (ELet ["_2"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "-"%string)) [(EVar "L"%string);(ELit (Integer (1)))]) (ELet ["_3"%string] (EApp (EFunId ("sublist_2"%string, 2)) [(EVar "T"%string);(EVar "_2"%string)]) (ECons (EVar "H"%string) (EVar "_3"%string)))));([(PVar "_8"%string);(PLit (Integer (0)))], (ELit (Atom "true"%string)), ENil);([(PVar "List"%string);(PVar "L"%string)], (ELet ["_4"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_list"%string)) [(EVar "List"%string)]) (ELet ["_5"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom ">"%string)) [(EVar "L"%string);(ELit (Integer (0)))]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "and"%string)) [(EVar "_4"%string);(EVar "_5"%string)]))), ENil);([(PVar "_7"%string);(PVar "_6"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_7"%string);(EVar "_6"%string)])]))]) |};
          {| identifier := ("delete"%string, 2) ; varl := ["_0"%string;"_1"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string)]) [([(PVar "Item"%string);(PCons (PVar "_5"%string) (PVar "Rest"%string))], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=:="%string)) [(EVar "_5"%string);(EVar "Item"%string)]), (EVar "Rest"%string));([(PVar "Item"%string);(PCons (PVar "H"%string) (PVar "Rest"%string))], (ELit (Atom "true"%string)), (ELet ["_2"%string] (EApp (EFunId ("delete"%string, 2)) [(EVar "Item"%string);(EVar "Rest"%string)]) (ECons (EVar "H"%string) (EVar "_2"%string))));([(PVar "_6"%string);PNil], (ELit (Atom "true"%string)), ENil);([(PVar "_4"%string);(PVar "_3"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_4"%string);(EVar "_3"%string)])]))]) |};
          {| identifier := ("zip"%string, 2) ; varl := ["_0"%string;"_1"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string)]) [([(PCons (PVar "X"%string) (PVar "Xs"%string));(PCons (PVar "Y"%string) (PVar "Ys"%string))], (ELit (Atom "true"%string)), (ELet ["_2"%string] (EApp (EFunId ("zip"%string, 2)) [(EVar "Xs"%string);(EVar "Ys"%string)]) (ECons (ETuple [(EVar "X"%string);(EVar "Y"%string)]) (EVar "_2"%string))));([PNil;PNil], (ELit (Atom "true"%string)), ENil);([(PVar "_4"%string);(PVar "_3"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_4"%string);(EVar "_3"%string)])]))]) |};
          {| identifier := ("unzip"%string, 1) ; varl := ["_0"%string]; body := (EApp (EFunId ("unzip"%string, 3)) [(EVar "_0"%string);ENil;ENil]) |};
          {| identifier := ("unzip"%string, 3) ; varl := ["_0"%string;"_1"%string;"_2"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string)]) [([(PCons (PTuple [(PVar "X"%string);(PVar "Y"%string)]) (PVar "Ts"%string));(PVar "Xs"%string);(PVar "Ys"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("unzip"%string, 3)) [(EVar "Ts"%string);(ECons (EVar "X"%string) (EVar "Xs"%string));(ECons (EVar "Y"%string) (EVar "Ys"%string))]));([PNil;(PVar "Xs"%string);(PVar "Ys"%string)], (ELit (Atom "true"%string)), (ELet ["_4"%string] (EApp (EFunId ("reverse"%string, 1)) [(EVar "Xs"%string)]) (ELet ["_3"%string] (EApp (EFunId ("reverse"%string, 1)) [(EVar "Ys"%string)]) (ETuple [(EVar "_4"%string);(EVar "_3"%string)]))));([(PVar "_7"%string);(PVar "_6"%string);(PVar "_5"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_7"%string);(EVar "_6"%string);(EVar "_5"%string)])]))]) |};
          {| identifier := ("zip3"%string, 3) ; varl := ["_0"%string;"_1"%string;"_2"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string)]) [([(PCons (PVar "X"%string) (PVar "Xs"%string));(PCons (PVar "Y"%string) (PVar "Ys"%string));(PCons (PVar "Z"%string) (PVar "Zs"%string))], (ELit (Atom "true"%string)), (ELet ["_3"%string] (EApp (EFunId ("zip3"%string, 3)) [(EVar "Xs"%string);(EVar "Ys"%string);(EVar "Zs"%string)]) (ECons (ETuple [(EVar "X"%string);(EVar "Y"%string);(EVar "Z"%string)]) (EVar "_3"%string))));([PNil;PNil;PNil], (ELit (Atom "true"%string)), ENil);([(PVar "_6"%string);(PVar "_5"%string);(PVar "_4"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_6"%string);(EVar "_5"%string);(EVar "_4"%string)])]))]) |};
          {| identifier := ("unzip3"%string, 1) ; varl := ["_0"%string]; body := (EApp (EFunId ("unzip3"%string, 4)) [(EVar "_0"%string);ENil;ENil;ENil]) |};
          {| identifier := ("unzip3"%string, 4) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string)]) [([(PCons (PTuple [(PVar "X"%string);(PVar "Y"%string);(PVar "Z"%string)]) (PVar "Ts"%string));(PVar "Xs"%string);(PVar "Ys"%string);(PVar "Zs"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("unzip3"%string, 4)) [(EVar "Ts"%string);(ECons (EVar "X"%string) (EVar "Xs"%string));(ECons (EVar "Y"%string) (EVar "Ys"%string));(ECons (EVar "Z"%string) (EVar "Zs"%string))]));([PNil;(PVar "Xs"%string);(PVar "Ys"%string);(PVar "Zs"%string)], (ELit (Atom "true"%string)), (ELet ["_6"%string] (EApp (EFunId ("reverse"%string, 1)) [(EVar "Xs"%string)]) (ELet ["_5"%string] (EApp (EFunId ("reverse"%string, 1)) [(EVar "Ys"%string)]) (ELet ["_4"%string] (EApp (EFunId ("reverse"%string, 1)) [(EVar "Zs"%string)]) (ETuple [(EVar "_6"%string);(EVar "_5"%string);(EVar "_4"%string)])))));([(PVar "_10"%string);(PVar "_9"%string);(PVar "_8"%string);(PVar "_7"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_10"%string);(EVar "_9"%string);(EVar "_8"%string);(EVar "_7"%string)])]))]) |};
          {| identifier := ("zipwith"%string, 3) ; varl := ["_0"%string;"_1"%string;"_2"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string)]) [([(PVar "F"%string);(PCons (PVar "X"%string) (PVar "Xs"%string));(PCons (PVar "Y"%string) (PVar "Ys"%string))], (ELit (Atom "true"%string)), (ELet ["_3"%string] (EApp (EVar "F"%string) [(EVar "X"%string);(EVar "Y"%string)]) (ELet ["_4"%string] (EApp (EFunId ("zipwith"%string, 3)) [(EVar "F"%string);(EVar "Xs"%string);(EVar "Ys"%string)]) (ECons (EVar "_3"%string) (EVar "_4"%string)))));([(PVar "F"%string);PNil;PNil], (ETry (ELet ["_5"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_function"%string)) [(EVar "F"%string);(ELit (Integer (2)))]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=:="%string)) [(EVar "_5"%string);(ELit (Atom "true"%string))])) ["Try"%string] (EVar "Try"%string) ["T"%string;"R"%string] (ELit (Atom "false"%string))), ENil);([(PVar "_8"%string);(PVar "_7"%string);(PVar "_6"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_8"%string);(EVar "_7"%string);(EVar "_6"%string)])]))]) |};
          {| identifier := ("zipwith3"%string, 4) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string)]) [([(PVar "F"%string);(PCons (PVar "X"%string) (PVar "Xs"%string));(PCons (PVar "Y"%string) (PVar "Ys"%string));(PCons (PVar "Z"%string) (PVar "Zs"%string))], (ELit (Atom "true"%string)), (ELet ["_4"%string] (EApp (EVar "F"%string) [(EVar "X"%string);(EVar "Y"%string);(EVar "Z"%string)]) (ELet ["_5"%string] (EApp (EFunId ("zipwith3"%string, 4)) [(EVar "F"%string);(EVar "Xs"%string);(EVar "Ys"%string);(EVar "Zs"%string)]) (ECons (EVar "_4"%string) (EVar "_5"%string)))));([(PVar "F"%string);PNil;PNil;PNil], (ETry (ELet ["_6"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_function"%string)) [(EVar "F"%string);(ELit (Integer (3)))]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=:="%string)) [(EVar "_6"%string);(ELit (Atom "true"%string))])) ["Try"%string] (EVar "Try"%string) ["T"%string;"R"%string] (ELit (Atom "false"%string))), ENil);([(PVar "_10"%string);(PVar "_9"%string);(PVar "_8"%string);(PVar "_7"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_10"%string);(EVar "_9"%string);(EVar "_8"%string);(EVar "_7"%string)])]))]) |};
          {| identifier := ("sort"%string, 1) ; varl := ["_0"%string]; body := (ECase (EVar "_0"%string) [([(PTuple [(PLit (Atom "c_alias"%string));PNil;(PVar "L0"%string);(PCons (PVar "X"%string) (PCons (PVar "Y"%string) (PVar "L"%string)))])], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "X"%string);(EVar "Y"%string)]), (ECase (EVar "L"%string) [([PNil], (ELit (Atom "true"%string)), (EVar "L0"%string));([(PCons (PVar "Z"%string) PNil)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "Y"%string);(EVar "Z"%string)]), (EVar "L0"%string));([(PCons (PVar "Z"%string) PNil)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "X"%string);(EVar "Z"%string)]), (ECons (EVar "X"%string) (ECons (EVar "Z"%string) (ECons (EVar "Y"%string) ENil))));([(PCons (PVar "Z"%string) PNil)], (ELit (Atom "true"%string)), (ECons (EVar "Z"%string) (ECons (EVar "X"%string) (ECons (EVar "Y"%string) ENil))));([(PVar "_4"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "X"%string);(EVar "Y"%string)]), (EApp (EFunId ("sort_1"%string, 3)) [(EVar "Y"%string);(EVar "L"%string);(ECons (EVar "X"%string) ENil)]));([(PVar "_5"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("split_1"%string, 5)) [(EVar "X"%string);(EVar "Y"%string);(EVar "L"%string);ENil;ENil]))]));([(PCons (PVar "X"%string) (PCons (PVar "Y"%string) (PVar "L"%string)))], (ELit (Atom "true"%string)), (ECase (EVar "L"%string) [([PNil], (ELit (Atom "true"%string)), (ECons (EVar "Y"%string) (ECons (EVar "X"%string) ENil)));([(PCons (PVar "Z"%string) PNil)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "X"%string);(EVar "Z"%string)]), (ECons (EVar "Y"%string) (ECons (EVar "X"%string) (EVar "L"%string))));([(PCons (PVar "Z"%string) PNil)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "Y"%string);(EVar "Z"%string)]), (ECons (EVar "Y"%string) (ECons (EVar "Z"%string) (ECons (EVar "X"%string) ENil))));([(PCons (PVar "Z"%string) PNil)], (ELit (Atom "true"%string)), (ECons (EVar "Z"%string) (ECons (EVar "Y"%string) (ECons (EVar "X"%string) ENil))));([(PVar "_6"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("split_2"%string, 5)) [(EVar "X"%string);(EVar "Y"%string);(EVar "L"%string);ENil;ENil]))]));([(PTuple [(PLit (Atom "c_alias"%string));PNil;(PVar "L"%string);(PCons (PVar "_7"%string) PNil)])], (ELit (Atom "true"%string)), (EVar "L"%string));([(PTuple [(PLit (Atom "c_alias"%string));PNil;(PVar "L"%string);PNil])], (ELit (Atom "true"%string)), (EVar "L"%string));([(PVar "_3"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_3"%string)])]))]) |};
          {| identifier := ("sort_1"%string, 3) ; varl := ["_0"%string;"_1"%string;"_2"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string)]) [([(PVar "X"%string);(PCons (PVar "Y"%string) (PVar "L"%string));(PVar "R"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "X"%string);(EVar "Y"%string)]), (EApp (EFunId ("sort_1"%string, 3)) [(EVar "Y"%string);(EVar "L"%string);(ECons (EVar "X"%string) (EVar "R"%string))]));([(PVar "X"%string);(PCons (PVar "Y"%string) (PVar "L"%string));(PVar "R"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "<"%string)) [(EVar "X"%string);(EVar "Y"%string)]), (EApp (EFunId ("split_1"%string, 5)) [(EVar "X"%string);(EVar "Y"%string);(EVar "L"%string);(EVar "R"%string);ENil]));([(PVar "X"%string);(PCons (PVar "Y"%string) (PVar "L"%string));(PVar "R"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("split_2"%string, 5)) [(EVar "X"%string);(EVar "Y"%string);(EVar "L"%string);(EVar "R"%string);ENil]));([(PVar "X"%string);PNil;(PVar "R"%string)], (ELit (Atom "true"%string)), (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "R"%string);(ECons (EVar "X"%string) ENil)]));([(PVar "_5"%string);(PVar "_4"%string);(PVar "_3"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_5"%string);(EVar "_4"%string);(EVar "_3"%string)])]))]) |};
          {| identifier := ("merge"%string, 1) ; varl := ["_0"%string]; body := (EApp (EFunId ("mergel"%string, 2)) [(EVar "_0"%string);ENil]) |};
          {| identifier := ("merge3"%string, 3) ; varl := ["_0"%string;"_1"%string;"_2"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string)]) [([(PVar "L1"%string);PNil;(PVar "L3"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("merge"%string, 2)) [(EVar "L1"%string);(EVar "L3"%string)]));([(PVar "L1"%string);(PVar "L2"%string);PNil], (ELit (Atom "true"%string)), (EApp (EFunId ("merge"%string, 2)) [(EVar "L1"%string);(EVar "L2"%string)]));([(PVar "L1"%string);(PCons (PVar "H2"%string) (PVar "T2"%string));(PCons (PVar "H3"%string) (PVar "T3"%string))], (ELit (Atom "true"%string)), (ELet ["_3"%string] (EApp (EFunId ("merge3_1"%string, 6)) [(EVar "L1"%string);ENil;(EVar "H2"%string);(EVar "T2"%string);(EVar "H3"%string);(EVar "T3"%string)]) (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "_3"%string);ENil])));([(PVar "_6"%string);(PVar "_5"%string);(PVar "_4"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_6"%string);(EVar "_5"%string);(EVar "_4"%string)])]))]) |};
          {| identifier := ("rmerge3"%string, 3) ; varl := ["_0"%string;"_1"%string;"_2"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string)]) [([(PVar "L1"%string);PNil;(PVar "L3"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rmerge"%string, 2)) [(EVar "L1"%string);(EVar "L3"%string)]));([(PVar "L1"%string);(PVar "L2"%string);PNil], (ELit (Atom "true"%string)), (EApp (EFunId ("rmerge"%string, 2)) [(EVar "L1"%string);(EVar "L2"%string)]));([(PVar "L1"%string);(PCons (PVar "H2"%string) (PVar "T2"%string));(PCons (PVar "H3"%string) (PVar "T3"%string))], (ELit (Atom "true"%string)), (ELet ["_3"%string] (EApp (EFunId ("rmerge3_1"%string, 6)) [(EVar "L1"%string);ENil;(EVar "H2"%string);(EVar "T2"%string);(EVar "H3"%string);(EVar "T3"%string)]) (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "_3"%string);ENil])));([(PVar "_6"%string);(PVar "_5"%string);(PVar "_4"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_6"%string);(EVar "_5"%string);(EVar "_4"%string)])]))]) |};
          {| identifier := ("merge"%string, 2) ; varl := ["_0"%string;"_1"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string)]) [([(PVar "T1"%string);PNil], (ELit (Atom "true"%string)), (EVar "T1"%string));([(PVar "T1"%string);(PCons (PVar "H2"%string) (PVar "T2"%string))], (ELit (Atom "true"%string)), (ELet ["_2"%string] (EApp (EFunId ("merge2_1"%string, 4)) [(EVar "T1"%string);(EVar "H2"%string);(EVar "T2"%string);ENil]) (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "_2"%string);ENil])));([(PVar "_4"%string);(PVar "_3"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_4"%string);(EVar "_3"%string)])]))]) |};
          {| identifier := ("rmerge"%string, 2) ; varl := ["_0"%string;"_1"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string)]) [([(PVar "T1"%string);PNil], (ELit (Atom "true"%string)), (EVar "T1"%string));([(PVar "T1"%string);(PCons (PVar "H2"%string) (PVar "T2"%string))], (ELit (Atom "true"%string)), (ELet ["_2"%string] (EApp (EFunId ("rmerge2_1"%string, 4)) [(EVar "T1"%string);(EVar "H2"%string);(EVar "T2"%string);ENil]) (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "_2"%string);ENil])));([(PVar "_4"%string);(PVar "_3"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_4"%string);(EVar "_3"%string)])]))]) |};
          {| identifier := ("concat"%string, 1) ; varl := ["_0"%string]; body := (ELet ["_1"%string] (EFunId ("thing_to_list"%string, 1)) (EApp (EFunId ("flatmap"%string, 2)) [(EVar "_1"%string);(EVar "_0"%string)])) |};
          {| identifier := ("thing_to_list"%string, 1) ; varl := ["_0"%string]; body := (ECase (EVar "_0"%string) [([(PVar "X"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_integer"%string)) [(EVar "_0"%string)]), (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "integer_to_list"%string)) [(EVar "X"%string)]));([(PVar "X"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_float"%string)) [(EVar "_0"%string)]), (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "float_to_list"%string)) [(EVar "X"%string)]));([(PVar "X"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_atom"%string)) [(EVar "_0"%string)]), (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "atom_to_list"%string)) [(EVar "X"%string)]));([(PVar "X"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_list"%string)) [(EVar "_0"%string)]), (EVar "X"%string));([(PVar "_1"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_1"%string)])]))]) |};
          {| identifier := ("flatten"%string, 1) ; varl := ["_0"%string]; body := (ECase (EVar "_0"%string) [([(PVar "List"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_list"%string)) [(EVar "_0"%string)]), (EApp (EFunId ("do_flatten"%string, 2)) [(EVar "List"%string);ENil]));([(PVar "_1"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_1"%string)])]))]) |};
          {| identifier := ("flatten"%string, 2) ; varl := ["_0"%string;"_1"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string)]) [([(PVar "List"%string);(PVar "Tail"%string)], (ELet ["_2"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_list"%string)) [(EVar "List"%string)]) (ELet ["_3"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_list"%string)) [(EVar "Tail"%string)]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "and"%string)) [(EVar "_2"%string);(EVar "_3"%string)]))), (EApp (EFunId ("do_flatten"%string, 2)) [(EVar "List"%string);(EVar "Tail"%string)]));([(PVar "_5"%string);(PVar "_4"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_5"%string);(EVar "_4"%string)])]))]) |};
          {| identifier := ("do_flatten"%string, 2) ; varl := ["_0"%string;"_1"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string)]) [([(PCons (PVar "H"%string) (PVar "T"%string));(PVar "Tail"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_list"%string)) [(EVar "H"%string)]), (ELet ["_2"%string] (EApp (EFunId ("do_flatten"%string, 2)) [(EVar "T"%string);(EVar "Tail"%string)]) (EApp (EFunId ("do_flatten"%string, 2)) [(EVar "H"%string);(EVar "_2"%string)])));([(PCons (PVar "H"%string) (PVar "T"%string));(PVar "Tail"%string)], (ELit (Atom "true"%string)), (ELet ["_3"%string] (EApp (EFunId ("do_flatten"%string, 2)) [(EVar "T"%string);(EVar "Tail"%string)]) (ECons (EVar "H"%string) (EVar "_3"%string))));([PNil;(PVar "Tail"%string)], (ELit (Atom "true"%string)), (EVar "Tail"%string));([(PVar "_5"%string);(PVar "_4"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_5"%string);(EVar "_4"%string)])]))]) |};
          {| identifier := ("flatlength"%string, 1) ; varl := ["_0"%string]; body := (EApp (EFunId ("flatlength"%string, 2)) [(EVar "_0"%string);(ELit (Integer (0)))]) |};
          {| identifier := ("flatlength"%string, 2) ; varl := ["_0"%string;"_1"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string)]) [([(PCons (PVar "H"%string) (PVar "T"%string));(PVar "L"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_list"%string)) [(EVar "H"%string)]), (ELet ["_2"%string] (EApp (EFunId ("flatlength"%string, 2)) [(EVar "T"%string);(EVar "L"%string)]) (EApp (EFunId ("flatlength"%string, 2)) [(EVar "H"%string);(EVar "_2"%string)])));([(PCons (PVar "_6"%string) (PVar "T"%string));(PVar "L"%string)], (ELit (Atom "true"%string)), (ELet ["_3"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "+"%string)) [(EVar "L"%string);(ELit (Integer (1)))]) (EApp (EFunId ("flatlength"%string, 2)) [(EVar "T"%string);(EVar "_3"%string)])));([PNil;(PVar "L"%string)], (ELit (Atom "true"%string)), (EVar "L"%string));([(PVar "_5"%string);(PVar "_4"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_5"%string);(EVar "_4"%string)])]))]) |};
          {| identifier := ("keydelete"%string, 3) ; varl := ["_0"%string;"_1"%string;"_2"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string)]) [([(PVar "K"%string);(PVar "N"%string);(PVar "L"%string)], (ELet ["_3"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_integer"%string)) [(EVar "N"%string)]) (ELet ["_4"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom ">"%string)) [(EVar "N"%string);(ELit (Integer (0)))]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "and"%string)) [(EVar "_3"%string);(EVar "_4"%string)]))), (EApp (EFunId ("keydelete3"%string, 3)) [(EVar "K"%string);(EVar "N"%string);(EVar "L"%string)]));([(PVar "_7"%string);(PVar "_6"%string);(PVar "_5"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_7"%string);(EVar "_6"%string);(EVar "_5"%string)])]))]) |};
          {| identifier := ("keydelete3"%string, 3) ; varl := ["_0"%string;"_1"%string;"_2"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string)]) [([(PVar "Key"%string);(PVar "N"%string);(PCons (PVar "H"%string) (PVar "T"%string))], (ETry (ELet ["_3"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "N"%string);(EVar "H"%string)]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "_3"%string);(EVar "Key"%string)])) ["Try"%string] (EVar "Try"%string) ["T"%string;"R"%string] (ELit (Atom "false"%string))), (EVar "T"%string));([(PVar "Key"%string);(PVar "N"%string);(PCons (PVar "H"%string) (PVar "T"%string))], (ELit (Atom "true"%string)), (ELet ["_4"%string] (EApp (EFunId ("keydelete3"%string, 3)) [(EVar "Key"%string);(EVar "N"%string);(EVar "T"%string)]) (ECons (EVar "H"%string) (EVar "_4"%string))));([(PVar "_8"%string);(PVar "_9"%string);PNil], (ELit (Atom "true"%string)), ENil);([(PVar "_7"%string);(PVar "_6"%string);(PVar "_5"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_7"%string);(EVar "_6"%string);(EVar "_5"%string)])]))]) |};
          {| identifier := ("keyreplace"%string, 4) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string)]) [([(PVar "K"%string);(PVar "N"%string);(PVar "L"%string);(PVar "New"%string)], (ETry (ELet ["_4"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_integer"%string)) [(EVar "N"%string)]) (ELet ["_5"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom ">"%string)) [(EVar "N"%string);(ELit (Integer (0)))]) (ELet ["_6"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_tuple"%string)) [(EVar "New"%string)]) (ELet ["_7"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "and"%string)) [(EVar "_5"%string);(EVar "_6"%string)]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "and"%string)) [(EVar "_4"%string);(EVar "_7"%string)]))))) ["Try"%string] (EVar "Try"%string) ["T"%string;"R"%string] (ELit (Atom "false"%string))), (EApp (EFunId ("keyreplace3"%string, 4)) [(EVar "K"%string);(EVar "N"%string);(EVar "L"%string);(EVar "New"%string)]));([(PVar "_11"%string);(PVar "_10"%string);(PVar "_9"%string);(PVar "_8"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_11"%string);(EVar "_10"%string);(EVar "_9"%string);(EVar "_8"%string)])]))]) |};
          {| identifier := ("keyreplace3"%string, 4) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string)]) [([(PVar "Key"%string);(PVar "Pos"%string);(PCons (PVar "Tup"%string) (PVar "Tail"%string));(PVar "New"%string)], (ETry (ELet ["_4"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "Pos"%string);(EVar "Tup"%string)]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "_4"%string);(EVar "Key"%string)])) ["Try"%string] (EVar "Try"%string) ["T"%string;"R"%string] (ELit (Atom "false"%string))), (ECons (EVar "New"%string) (EVar "Tail"%string)));([(PVar "Key"%string);(PVar "Pos"%string);(PCons (PVar "H"%string) (PVar "T"%string));(PVar "New"%string)], (ELit (Atom "true"%string)), (ELet ["_5"%string] (EApp (EFunId ("keyreplace3"%string, 4)) [(EVar "Key"%string);(EVar "Pos"%string);(EVar "T"%string);(EVar "New"%string)]) (ECons (EVar "H"%string) (EVar "_5"%string))));([(PVar "_10"%string);(PVar "_11"%string);PNil;(PVar "_12"%string)], (ELit (Atom "true"%string)), ENil);([(PVar "_9"%string);(PVar "_8"%string);(PVar "_7"%string);(PVar "_6"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_9"%string);(EVar "_8"%string);(EVar "_7"%string);(EVar "_6"%string)])]))]) |};
          {| identifier := ("keytake"%string, 3) ; varl := ["_0"%string;"_1"%string;"_2"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string)]) [([(PVar "Key"%string);(PVar "N"%string);(PVar "L"%string)], (ELet ["_3"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_integer"%string)) [(EVar "N"%string)]) (ELet ["_4"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom ">"%string)) [(EVar "N"%string);(ELit (Integer (0)))]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "and"%string)) [(EVar "_3"%string);(EVar "_4"%string)]))), (EApp (EFunId ("keytake"%string, 4)) [(EVar "Key"%string);(EVar "N"%string);(EVar "L"%string);ENil]));([(PVar "_7"%string);(PVar "_6"%string);(PVar "_5"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_7"%string);(EVar "_6"%string);(EVar "_5"%string)])]))]) |};
          {| identifier := ("keytake"%string, 4) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string)]) [([(PVar "Key"%string);(PVar "N"%string);(PCons (PVar "H"%string) (PVar "T"%string));(PVar "L"%string)], (ETry (ELet ["_4"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "N"%string);(EVar "H"%string)]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "_4"%string);(EVar "Key"%string)])) ["Try"%string] (EVar "Try"%string) ["T"%string;"R"%string] (ELit (Atom "false"%string))), (ELet ["_5"%string] (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "L"%string);(EVar "T"%string)]) (ETuple [(ELit (Atom "value"%string));(EVar "H"%string);(EVar "_5"%string)])));([(PVar "Key"%string);(PVar "N"%string);(PCons (PVar "H"%string) (PVar "T"%string));(PVar "L"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("keytake"%string, 4)) [(EVar "Key"%string);(EVar "N"%string);(EVar "T"%string);(ECons (EVar "H"%string) (EVar "L"%string))]));([(PVar "_K"%string);(PVar "_N"%string);PNil;(PVar "_L"%string)], (ELit (Atom "true"%string)), (ELit (Atom "false"%string)));([(PVar "_9"%string);(PVar "_8"%string);(PVar "_7"%string);(PVar "_6"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_9"%string);(EVar "_8"%string);(EVar "_7"%string);(EVar "_6"%string)])]))]) |};
          {| identifier := ("keystore"%string, 4) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string)]) [([(PVar "K"%string);(PVar "N"%string);(PVar "L"%string);(PVar "New"%string)], (ETry (ELet ["_4"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_integer"%string)) [(EVar "N"%string)]) (ELet ["_5"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom ">"%string)) [(EVar "N"%string);(ELit (Integer (0)))]) (ELet ["_6"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_tuple"%string)) [(EVar "New"%string)]) (ELet ["_7"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "and"%string)) [(EVar "_5"%string);(EVar "_6"%string)]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "and"%string)) [(EVar "_4"%string);(EVar "_7"%string)]))))) ["Try"%string] (EVar "Try"%string) ["T"%string;"R"%string] (ELit (Atom "false"%string))), (EApp (EFunId ("keystore2"%string, 4)) [(EVar "K"%string);(EVar "N"%string);(EVar "L"%string);(EVar "New"%string)]));([(PVar "_11"%string);(PVar "_10"%string);(PVar "_9"%string);(PVar "_8"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_11"%string);(EVar "_10"%string);(EVar "_9"%string);(EVar "_8"%string)])]))]) |};
          {| identifier := ("keystore2"%string, 4) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string)]) [([(PVar "Key"%string);(PVar "N"%string);(PCons (PVar "H"%string) (PVar "T"%string));(PVar "New"%string)], (ETry (ELet ["_4"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "N"%string);(EVar "H"%string)]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "_4"%string);(EVar "Key"%string)])) ["Try"%string] (EVar "Try"%string) ["T"%string;"R"%string] (ELit (Atom "false"%string))), (ECons (EVar "New"%string) (EVar "T"%string)));([(PVar "Key"%string);(PVar "N"%string);(PCons (PVar "H"%string) (PVar "T"%string));(PVar "New"%string)], (ELit (Atom "true"%string)), (ELet ["_5"%string] (EApp (EFunId ("keystore2"%string, 4)) [(EVar "Key"%string);(EVar "N"%string);(EVar "T"%string);(EVar "New"%string)]) (ECons (EVar "H"%string) (EVar "_5"%string))));([(PVar "_Key"%string);(PVar "_N"%string);PNil;(PVar "New"%string)], (ELit (Atom "true"%string)), (ECons (EVar "New"%string) ENil));([(PVar "_9"%string);(PVar "_8"%string);(PVar "_7"%string);(PVar "_6"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_9"%string);(EVar "_8"%string);(EVar "_7"%string);(EVar "_6"%string)])]))]) |};
          {| identifier := ("keysort"%string, 2) ; varl := ["_0"%string;"_1"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string)]) [([(PVar "I"%string);(PVar "L"%string)], (ELet ["_2"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_integer"%string)) [(EVar "I"%string)]) (ELet ["_3"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom ">"%string)) [(EVar "I"%string);(ELit (Integer (0)))]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "and"%string)) [(EVar "_2"%string);(EVar "_3"%string)]))), (ECase (EVar "L"%string) [([PNil], (ELit (Atom "true"%string)), (EVar "L"%string));([(PCons (PVar "_14"%string) PNil)], (ELit (Atom "true"%string)), (EVar "L"%string));([(PCons (PVar "X"%string) (PCons (PVar "Y"%string) (PVar "T"%string)))], (ELit (Atom "true"%string)), (ELet ["_5"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "I"%string);(EVar "X"%string)]) (ELet ["_4"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "I"%string);(EVar "Y"%string)]) (ECase (EValues [(EVar "_5"%string);(EVar "_4"%string)]) [([(PVar "EX"%string);(PVar "EY"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "EX"%string);(EVar "EY"%string)]), (ECase (EVar "T"%string) [([PNil], (ELit (Atom "true"%string)), (EVar "L"%string));([(PCons (PVar "Z"%string) PNil)], (ELit (Atom "true"%string)), (ECase (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "I"%string);(EVar "Z"%string)]) [([(PVar "EZ"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "EY"%string);(EVar "EZ"%string)]), (EVar "L"%string));([(PVar "EZ"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "EX"%string);(EVar "EZ"%string)]), (ECons (EVar "X"%string) (ECons (EVar "Z"%string) (ECons (EVar "Y"%string) ENil))));([(PVar "_EZ"%string)], (ELit (Atom "true"%string)), (ECons (EVar "Z"%string) (ECons (EVar "X"%string) (ECons (EVar "Y"%string) ENil))))]));([(PVar "_15"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "X"%string);(EVar "Y"%string)]), (EApp (EFunId ("keysort_1"%string, 5)) [(EVar "I"%string);(EVar "Y"%string);(EVar "EY"%string);(EVar "T"%string);(ECons (EVar "X"%string) ENil)]));([(PVar "_16"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("keysplit_1"%string, 8)) [(EVar "I"%string);(EVar "X"%string);(EVar "EX"%string);(EVar "Y"%string);(EVar "EY"%string);(EVar "T"%string);ENil;ENil]))]));([(PVar "EX"%string);(PVar "EY"%string)], (ELit (Atom "true"%string)), (ECase (EVar "T"%string) [([PNil], (ELit (Atom "true"%string)), (ECons (EVar "Y"%string) (ECons (EVar "X"%string) ENil)));([(PCons (PVar "Z"%string) PNil)], (ELit (Atom "true"%string)), (ECase (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "I"%string);(EVar "Z"%string)]) [([(PVar "EZ"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "EX"%string);(EVar "EZ"%string)]), (ECons (EVar "Y"%string) (ECons (EVar "X"%string) (EVar "T"%string))));([(PVar "EZ"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "EY"%string);(EVar "EZ"%string)]), (ECons (EVar "Y"%string) (ECons (EVar "Z"%string) (ECons (EVar "X"%string) ENil))));([(PVar "_EZ"%string)], (ELit (Atom "true"%string)), (ECons (EVar "Z"%string) (ECons (EVar "Y"%string) (ECons (EVar "X"%string) ENil))))]));([(PVar "_17"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("keysplit_2"%string, 8)) [(EVar "I"%string);(EVar "X"%string);(EVar "EX"%string);(EVar "Y"%string);(EVar "EY"%string);(EVar "T"%string);ENil;ENil]))]))]))));([(PVar "_11"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "case_clause"%string));(EVar "_11"%string)])]))]));([(PVar "_13"%string);(PVar "_12"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_13"%string);(EVar "_12"%string)])]))]) |};
          {| identifier := ("keysort_1"%string, 5) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string)]) [([(PVar "I"%string);(PVar "X"%string);(PVar "EX"%string);(PCons (PVar "Y"%string) (PVar "L"%string));(PVar "R"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "X"%string);(EVar "Y"%string)]), (EApp (EFunId ("keysort_1"%string, 5)) [(EVar "I"%string);(EVar "Y"%string);(EVar "EX"%string);(EVar "L"%string);(ECons (EVar "X"%string) (EVar "R"%string))]));([(PVar "I"%string);(PVar "X"%string);(PVar "EX"%string);(PCons (PVar "Y"%string) (PVar "L"%string));(PVar "R"%string)], (ELit (Atom "true"%string)), (ECase (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "I"%string);(EVar "Y"%string)]) [([(PVar "EY"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "EX"%string);(EVar "EY"%string)]), (EApp (EFunId ("keysplit_1"%string, 8)) [(EVar "I"%string);(EVar "X"%string);(EVar "EX"%string);(EVar "Y"%string);(EVar "EY"%string);(EVar "L"%string);(EVar "R"%string);ENil]));([(PVar "EY"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("keysplit_2"%string, 8)) [(EVar "I"%string);(EVar "X"%string);(EVar "EX"%string);(EVar "Y"%string);(EVar "EY"%string);(EVar "L"%string);(EVar "R"%string);ENil]))]));([(PVar "_I"%string);(PVar "X"%string);(PVar "_EX"%string);PNil;(PVar "R"%string)], (ELit (Atom "true"%string)), (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "R"%string);(ECons (EVar "X"%string) ENil)]));([(PVar "_10"%string);(PVar "_9"%string);(PVar "_8"%string);(PVar "_7"%string);(PVar "_6"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_10"%string);(EVar "_9"%string);(EVar "_8"%string);(EVar "_7"%string);(EVar "_6"%string)])]))]) |};
          {| identifier := ("keymerge"%string, 3) ; varl := ["_0"%string;"_1"%string;"_2"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string)]) [([(PVar "Index"%string);(PVar "T1"%string);(PVar "L2"%string)], (ELet ["_3"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_integer"%string)) [(EVar "Index"%string)]) (ELet ["_4"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom ">"%string)) [(EVar "Index"%string);(ELit (Integer (0)))]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "and"%string)) [(EVar "_3"%string);(EVar "_4"%string)]))), (ECase (EVar "L2"%string) [([PNil], (ELit (Atom "true"%string)), (EVar "T1"%string));([(PCons (PVar "H2"%string) (PVar "T2"%string))], (ELit (Atom "true"%string)), (ELet ["E2"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "Index"%string);(EVar "H2"%string)]) (ELet ["M"%string] (EApp (EFunId ("keymerge2_1"%string, 6)) [(EVar "Index"%string);(EVar "T1"%string);(EVar "E2"%string);(EVar "H2"%string);(EVar "T2"%string);ENil]) (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "M"%string);ENil]))));([(PVar "_7"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "case_clause"%string));(EVar "_7"%string)])]))]));([(PVar "_10"%string);(PVar "_9"%string);(PVar "_8"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_10"%string);(EVar "_9"%string);(EVar "_8"%string)])]))]) |};
          {| identifier := ("rkeymerge"%string, 3) ; varl := ["_0"%string;"_1"%string;"_2"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string)]) [([(PVar "Index"%string);(PVar "T1"%string);(PVar "L2"%string)], (ELet ["_3"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_integer"%string)) [(EVar "Index"%string)]) (ELet ["_4"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom ">"%string)) [(EVar "Index"%string);(ELit (Integer (0)))]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "and"%string)) [(EVar "_3"%string);(EVar "_4"%string)]))), (ECase (EVar "L2"%string) [([PNil], (ELit (Atom "true"%string)), (EVar "T1"%string));([(PCons (PVar "H2"%string) (PVar "T2"%string))], (ELit (Atom "true"%string)), (ELet ["E2"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "Index"%string);(EVar "H2"%string)]) (ELet ["M"%string] (EApp (EFunId ("rkeymerge2_1"%string, 6)) [(EVar "Index"%string);(EVar "T1"%string);(EVar "E2"%string);(EVar "H2"%string);(EVar "T2"%string);ENil]) (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "M"%string);ENil]))));([(PVar "_7"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "case_clause"%string));(EVar "_7"%string)])]))]));([(PVar "_10"%string);(PVar "_9"%string);(PVar "_8"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_10"%string);(EVar "_9"%string);(EVar "_8"%string)])]))]) |};
          {| identifier := ("ukeysort"%string, 2) ; varl := ["_0"%string;"_1"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string)]) [([(PVar "I"%string);(PVar "L"%string)], (ELet ["_2"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_integer"%string)) [(EVar "I"%string)]) (ELet ["_3"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom ">"%string)) [(EVar "I"%string);(ELit (Integer (0)))]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "and"%string)) [(EVar "_2"%string);(EVar "_3"%string)]))), (ECase (EVar "L"%string) [([PNil], (ELit (Atom "true"%string)), (EVar "L"%string));([(PCons (PVar "_14"%string) PNil)], (ELit (Atom "true"%string)), (EVar "L"%string));([(PCons (PVar "X"%string) (PCons (PVar "Y"%string) (PVar "T"%string)))], (ELit (Atom "true"%string)), (ELet ["_5"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "I"%string);(EVar "X"%string)]) (ELet ["_4"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "I"%string);(EVar "Y"%string)]) (ECase (EValues [(EVar "_5"%string);(EVar "_4"%string)]) [([(PVar "EX"%string);(PVar "EY"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "EX"%string);(EVar "EY"%string)]), (EApp (EFunId ("ukeysort_1"%string, 4)) [(EVar "I"%string);(EVar "X"%string);(EVar "EX"%string);(EVar "T"%string)]));([(PVar "EX"%string);(PVar "EY"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "<"%string)) [(EVar "EX"%string);(EVar "EY"%string)]), (ECase (EVar "T"%string) [([PNil], (ELit (Atom "true"%string)), (EVar "L"%string));([(PTuple [(PLit (Atom "c_alias"%string));(PCons (PTuple [(PLit (Integer (891)));(PLit (Integer (25)))]) (PCons (PTuple [(PLit (Atom "file"%string));(PCons (PLit (Integer (47))) (PCons (PLit (Integer (85))) (PCons (PLit (Integer (115))) (PCons (PLit (Integer (101))) (PCons (PLit (Integer (114))) (PCons (PLit (Integer (115))) (PCons (PLit (Integer (47))) (PCons (PLit (Integer (103))) (PCons (PLit (Integer (121))) (PCons (PLit (Integer (117))) (PCons (PLit (Integer (114))) (PCons (PLit (Integer (105))) (PCons (PLit (Integer (47))) (PCons (PLit (Integer (68))) (PCons (PLit (Integer (111))) (PCons (PLit (Integer (99))) (PCons (PLit (Integer (117))) (PCons (PLit (Integer (109))) (PCons (PLit (Integer (101))) (PCons (PLit (Integer (110))) (PCons (PLit (Integer (116))) (PCons (PLit (Integer (115))) (PCons (PLit (Integer (47))) (PCons (PLit (Integer (111))) (PCons (PLit (Integer (115))) (PCons (PLit (Integer (107))) (PCons (PLit (Integer (111))) (PCons (PLit (Integer (108))) (PCons (PLit (Integer (97))) (PCons (PLit (Integer (47))) (PCons (PLit (Integer (72))) (PCons (PLit (Integer (65))) (PCons (PLit (Integer (82))) (PCons (PLit (Integer (80))) (PCons (PLit (Integer (47))) (PCons (PLit (Integer (111))) (PCons (PLit (Integer (116))) (PCons (PLit (Integer (112))) (PCons (PLit (Integer (45))) (PCons (PLit (Integer (109))) (PCons (PLit (Integer (97))) (PCons (PLit (Integer (115))) (PCons (PLit (Integer (116))) (PCons (PLit (Integer (101))) (PCons (PLit (Integer (114))) (PCons (PLit (Integer (47))) (PCons (PLit (Integer (108))) (PCons (PLit (Integer (105))) (PCons (PLit (Integer (98))) (PCons (PLit (Integer (47))) (PCons (PLit (Integer (115))) (PCons (PLit (Integer (116))) (PCons (PLit (Integer (100))) (PCons (PLit (Integer (108))) (PCons (PLit (Integer (105))) (PCons (PLit (Integer (98))) (PCons (PLit (Integer (47))) (PCons (PLit (Integer (115))) (PCons (PLit (Integer (114))) (PCons (PLit (Integer (99))) (PCons (PLit (Integer (47))) (PCons (PLit (Integer (108))) (PCons (PLit (Integer (105))) (PCons (PLit (Integer (115))) (PCons (PLit (Integer (116))) (PCons (PLit (Integer (115))) (PCons (PLit (Integer (46))) (PCons (PLit (Integer (101))) (PCons (PLit (Integer (114))) (PCons (PLit (Integer (108))) PNil))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))]) PNil));(PVar "@r0"%string);(PCons (PVar "Z"%string) PNil)])], (ELit (Atom "true"%string)), (ECase (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "I"%string);(EVar "Z"%string)]) [([(PVar "EZ"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "EY"%string);(EVar "EZ"%string)]), (ECons (EVar "X"%string) (ECons (EVar "Y"%string) ENil)));([(PVar "EZ"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "<"%string)) [(EVar "EY"%string);(EVar "EZ"%string)]), (ECons (EVar "X"%string) (ECons (EVar "Y"%string) (EVar "@r0"%string))));([(PVar "EZ"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "EZ"%string);(EVar "EX"%string)]), (ECons (EVar "X"%string) (ECons (EVar "Y"%string) ENil)));([(PVar "EZ"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "EX"%string);(EVar "EZ"%string)]), (ECons (EVar "X"%string) (ECons (EVar "Z"%string) (ECons (EVar "Y"%string) ENil))));([(PVar "_EZ"%string)], (ELit (Atom "true"%string)), (ECons (EVar "Z"%string) (ECons (EVar "X"%string) (ECons (EVar "Y"%string) ENil))))]));([(PVar "_15"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("ukeysplit_1"%string, 8)) [(EVar "I"%string);(EVar "X"%string);(EVar "EX"%string);(EVar "Y"%string);(EVar "EY"%string);(EVar "T"%string);ENil;ENil]))]));([(PVar "EX"%string);(PVar "EY"%string)], (ELit (Atom "true"%string)), (ECase (EVar "T"%string) [([PNil], (ELit (Atom "true"%string)), (ECons (EVar "Y"%string) (ECons (EVar "X"%string) ENil)));([(PTuple [(PLit (Atom "c_alias"%string));(PCons (PTuple [(PLit (Integer (911)));(PLit (Integer (25)))]) (PCons (PTuple [(PLit (Atom "file"%string));(PCons (PLit (Integer (47))) (PCons (PLit (Integer (85))) (PCons (PLit (Integer (115))) (PCons (PLit (Integer (101))) (PCons (PLit (Integer (114))) (PCons (PLit (Integer (115))) (PCons (PLit (Integer (47))) (PCons (PLit (Integer (103))) (PCons (PLit (Integer (121))) (PCons (PLit (Integer (117))) (PCons (PLit (Integer (114))) (PCons (PLit (Integer (105))) (PCons (PLit (Integer (47))) (PCons (PLit (Integer (68))) (PCons (PLit (Integer (111))) (PCons (PLit (Integer (99))) (PCons (PLit (Integer (117))) (PCons (PLit (Integer (109))) (PCons (PLit (Integer (101))) (PCons (PLit (Integer (110))) (PCons (PLit (Integer (116))) (PCons (PLit (Integer (115))) (PCons (PLit (Integer (47))) (PCons (PLit (Integer (111))) (PCons (PLit (Integer (115))) (PCons (PLit (Integer (107))) (PCons (PLit (Integer (111))) (PCons (PLit (Integer (108))) (PCons (PLit (Integer (97))) (PCons (PLit (Integer (47))) (PCons (PLit (Integer (72))) (PCons (PLit (Integer (65))) (PCons (PLit (Integer (82))) (PCons (PLit (Integer (80))) (PCons (PLit (Integer (47))) (PCons (PLit (Integer (111))) (PCons (PLit (Integer (116))) (PCons (PLit (Integer (112))) (PCons (PLit (Integer (45))) (PCons (PLit (Integer (109))) (PCons (PLit (Integer (97))) (PCons (PLit (Integer (115))) (PCons (PLit (Integer (116))) (PCons (PLit (Integer (101))) (PCons (PLit (Integer (114))) (PCons (PLit (Integer (47))) (PCons (PLit (Integer (108))) (PCons (PLit (Integer (105))) (PCons (PLit (Integer (98))) (PCons (PLit (Integer (47))) (PCons (PLit (Integer (115))) (PCons (PLit (Integer (116))) (PCons (PLit (Integer (100))) (PCons (PLit (Integer (108))) (PCons (PLit (Integer (105))) (PCons (PLit (Integer (98))) (PCons (PLit (Integer (47))) (PCons (PLit (Integer (115))) (PCons (PLit (Integer (114))) (PCons (PLit (Integer (99))) (PCons (PLit (Integer (47))) (PCons (PLit (Integer (108))) (PCons (PLit (Integer (105))) (PCons (PLit (Integer (115))) (PCons (PLit (Integer (116))) (PCons (PLit (Integer (115))) (PCons (PLit (Integer (46))) (PCons (PLit (Integer (101))) (PCons (PLit (Integer (114))) (PCons (PLit (Integer (108))) PNil))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))]) PNil));(PVar "@r1"%string);(PCons (PVar "Z"%string) PNil)])], (ELit (Atom "true"%string)), (ECase (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "I"%string);(EVar "Z"%string)]) [([(PVar "EZ"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "EX"%string);(EVar "EZ"%string)]), (ECons (EVar "Y"%string) (ECons (EVar "X"%string) ENil)));([(PVar "EZ"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "<"%string)) [(EVar "EX"%string);(EVar "EZ"%string)]), (ECons (EVar "Y"%string) (ECons (EVar "X"%string) (EVar "@r1"%string))));([(PVar "EZ"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "EY"%string);(EVar "EZ"%string)]), (ECons (EVar "Y"%string) (ECons (EVar "X"%string) ENil)));([(PVar "EZ"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "EY"%string);(EVar "EZ"%string)]), (ECons (EVar "Y"%string) (ECons (EVar "Z"%string) (ECons (EVar "X"%string) ENil))));([(PVar "_EZ"%string)], (ELit (Atom "true"%string)), (ECons (EVar "Z"%string) (ECons (EVar "Y"%string) (ECons (EVar "X"%string) ENil))))]));([(PVar "_16"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("ukeysplit_2"%string, 5)) [(EVar "I"%string);(EVar "Y"%string);(EVar "EY"%string);(EVar "T"%string);(ECons (EVar "X"%string) ENil)]))]))]))));([(PVar "_11"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "case_clause"%string));(EVar "_11"%string)])]))]));([(PVar "_13"%string);(PVar "_12"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_13"%string);(EVar "_12"%string)])]))]) |};
          {| identifier := ("ukeysort_1"%string, 4) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string)]) [([(PVar "I"%string);(PVar "X"%string);(PVar "EX"%string);(PCons (PVar "Y"%string) (PVar "L"%string))], (ELit (Atom "true"%string)), (ECase (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "I"%string);(EVar "Y"%string)]) [([(PVar "EY"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "EX"%string);(EVar "EY"%string)]), (EApp (EFunId ("ukeysort_1"%string, 4)) [(EVar "I"%string);(EVar "X"%string);(EVar "EX"%string);(EVar "L"%string)]));([(PVar "EY"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "<"%string)) [(EVar "EX"%string);(EVar "EY"%string)]), (EApp (EFunId ("ukeysplit_1"%string, 8)) [(EVar "I"%string);(EVar "X"%string);(EVar "EX"%string);(EVar "Y"%string);(EVar "EY"%string);(EVar "L"%string);ENil;ENil]));([(PVar "EY"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("ukeysplit_2"%string, 5)) [(EVar "I"%string);(EVar "Y"%string);(EVar "EY"%string);(EVar "L"%string);(ECons (EVar "X"%string) ENil)]))]));([(PVar "_I"%string);(PVar "X"%string);(PVar "_EX"%string);PNil], (ELit (Atom "true"%string)), (ECons (EVar "X"%string) ENil));([(PVar "_8"%string);(PVar "_7"%string);(PVar "_6"%string);(PVar "_5"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_8"%string);(EVar "_7"%string);(EVar "_6"%string);(EVar "_5"%string)])]))]) |};
          {| identifier := ("ukeymerge"%string, 3) ; varl := ["_0"%string;"_1"%string;"_2"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string)]) [([(PVar "Index"%string);(PVar "L1"%string);(PVar "T2"%string)], (ELet ["_3"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_integer"%string)) [(EVar "Index"%string)]) (ELet ["_4"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom ">"%string)) [(EVar "Index"%string);(ELit (Integer (0)))]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "and"%string)) [(EVar "_3"%string);(EVar "_4"%string)]))), (ECase (EVar "L1"%string) [([PNil], (ELit (Atom "true"%string)), (EVar "T2"%string));([(PCons (PVar "H1"%string) (PVar "T1"%string))], (ELit (Atom "true"%string)), (ELet ["E1"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "Index"%string);(EVar "H1"%string)]) (ELet ["M"%string] (EApp (EFunId ("ukeymerge2_2"%string, 6)) [(EVar "Index"%string);(EVar "T1"%string);(EVar "E1"%string);(EVar "H1"%string);(EVar "T2"%string);ENil]) (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "M"%string);ENil]))));([(PVar "_7"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "case_clause"%string));(EVar "_7"%string)])]))]));([(PVar "_10"%string);(PVar "_9"%string);(PVar "_8"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_10"%string);(EVar "_9"%string);(EVar "_8"%string)])]))]) |};
          {| identifier := ("rukeymerge"%string, 3) ; varl := ["_0"%string;"_1"%string;"_2"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string)]) [([(PVar "Index"%string);(PVar "T1"%string);(PVar "L2"%string)], (ELet ["_3"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_integer"%string)) [(EVar "Index"%string)]) (ELet ["_4"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom ">"%string)) [(EVar "Index"%string);(ELit (Integer (0)))]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "and"%string)) [(EVar "_3"%string);(EVar "_4"%string)]))), (ECase (EVar "L2"%string) [([PNil], (ELit (Atom "true"%string)), (EVar "T1"%string));([(PCons (PVar "H2"%string) (PVar "T2"%string))], (ELit (Atom "true"%string)), (ELet ["E2"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "Index"%string);(EVar "H2"%string)]) (ELet ["M"%string] (EApp (EFunId ("rukeymerge2_1"%string, 6)) [(EVar "Index"%string);(EVar "T1"%string);(EVar "E2"%string);(EVar "T2"%string);ENil;(EVar "H2"%string)]) (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "M"%string);ENil]))));([(PVar "_7"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "case_clause"%string));(EVar "_7"%string)])]))]));([(PVar "_10"%string);(PVar "_9"%string);(PVar "_8"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_10"%string);(EVar "_9"%string);(EVar "_8"%string)])]))]) |};
          {| identifier := ("keymap"%string, 3) ; varl := ["_0"%string;"_1"%string;"_2"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string)]) [([(PVar "Fun"%string);(PVar "Index"%string);(PCons (PVar "Tup"%string) (PVar "Tail"%string))], (ELit (Atom "true"%string)), (ELet ["_3"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "Index"%string);(EVar "Tup"%string)]) (ELet ["_4"%string] (EApp (EVar "Fun"%string) [(EVar "_3"%string)]) (ELet ["_5"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "setelement"%string)) [(EVar "Index"%string);(EVar "Tup"%string);(EVar "_4"%string)]) (ELet ["_6"%string] (EApp (EFunId ("keymap"%string, 3)) [(EVar "Fun"%string);(EVar "Index"%string);(EVar "Tail"%string)]) (ECons (EVar "_5"%string) (EVar "_6"%string)))))));([(PVar "Fun"%string);(PVar "Index"%string);PNil], (ETry (ELet ["_7"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_integer"%string)) [(EVar "Index"%string)]) (ELet ["_8"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom ">="%string)) [(EVar "Index"%string);(ELit (Integer (1)))]) (ELet ["_9"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_function"%string)) [(EVar "Fun"%string);(ELit (Integer (1)))]) (ELet ["_10"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=:="%string)) [(EVar "_9"%string);(ELit (Atom "true"%string))]) (ELet ["_11"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "and"%string)) [(EVar "_8"%string);(EVar "_10"%string)]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "and"%string)) [(EVar "_7"%string);(EVar "_11"%string)])))))) ["Try"%string] (EVar "Try"%string) ["T"%string;"R"%string] (ELit (Atom "false"%string))), ENil);([(PVar "_14"%string);(PVar "_13"%string);(PVar "_12"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_14"%string);(EVar "_13"%string);(EVar "_12"%string)])]))]) |};
          {| identifier := ("enumerate"%string, 1) ; varl := ["_0"%string]; body := (ECase (EVar "_0"%string) [([(PVar "List1"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_list"%string)) [(EVar "_0"%string)]), (EApp (EFunId ("enumerate_1"%string, 2)) [(ELit (Integer (1)));(EVar "List1"%string)]));([(PVar "_1"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_1"%string)])]))]) |};
          {| identifier := ("enumerate"%string, 2) ; varl := ["_0"%string;"_1"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string)]) [([(PVar "Index"%string);(PVar "List1"%string)], (ELet ["_2"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_integer"%string)) [(EVar "Index"%string)]) (ELet ["_3"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_list"%string)) [(EVar "List1"%string)]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "and"%string)) [(EVar "_2"%string);(EVar "_3"%string)]))), (EApp (EFunId ("enumerate_1"%string, 2)) [(EVar "Index"%string);(EVar "List1"%string)]));([(PVar "_5"%string);(PVar "_4"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_5"%string);(EVar "_4"%string)])]))]) |};
          {| identifier := ("enumerate_1"%string, 2) ; varl := ["_0"%string;"_1"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string)]) [([(PVar "Index"%string);(PCons (PVar "H"%string) (PVar "T"%string))], (ELit (Atom "true"%string)), (ELet ["_2"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "+"%string)) [(EVar "Index"%string);(ELit (Integer (1)))]) (ELet ["_3"%string] (EApp (EFunId ("enumerate_1"%string, 2)) [(EVar "_2"%string);(EVar "T"%string)]) (ECons (ETuple [(EVar "Index"%string);(EVar "H"%string)]) (EVar "_3"%string)))));([(PVar "_Index"%string);PNil], (ELit (Atom "true"%string)), ENil);([(PVar "_5"%string);(PVar "_4"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_5"%string);(EVar "_4"%string)])]))]) |};
          {| identifier := ("sort"%string, 2) ; varl := ["_0"%string;"_1"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string)]) [([(PVar "Fun"%string);PNil], (ETry (ELet ["_2"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_function"%string)) [(EVar "Fun"%string);(ELit (Integer (2)))]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=:="%string)) [(EVar "_2"%string);(ELit (Atom "true"%string))])) ["Try"%string] (EVar "Try"%string) ["T"%string;"R"%string] (ELit (Atom "false"%string))), ENil);([(PVar "Fun"%string);(PTuple [(PLit (Atom "c_alias"%string));PNil;(PVar "L"%string);(PCons (PVar "_7"%string) PNil)])], (ETry (ELet ["_3"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_function"%string)) [(EVar "Fun"%string);(ELit (Integer (2)))]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=:="%string)) [(EVar "_3"%string);(ELit (Atom "true"%string))])) ["Try"%string] (EVar "Try"%string) ["T"%string;"R"%string] (ELit (Atom "false"%string))), (EVar "L"%string));([(PVar "Fun"%string);(PCons (PVar "X"%string) (PCons (PVar "Y"%string) (PVar "T"%string)))], (ELit (Atom "true"%string)), (ECase (EApp (EVar "Fun"%string) [(EVar "X"%string);(EVar "Y"%string)]) [([(PLit (Atom "true"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("fsplit_1"%string, 6)) [(EVar "Y"%string);(EVar "X"%string);(EVar "Fun"%string);(EVar "T"%string);ENil;ENil]));([(PLit (Atom "false"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("fsplit_2"%string, 6)) [(EVar "Y"%string);(EVar "X"%string);(EVar "Fun"%string);(EVar "T"%string);ENil;ENil]));([(PVar "_4"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "case_clause"%string));(EVar "_4"%string)])]))]));([(PVar "_6"%string);(PVar "_5"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_6"%string);(EVar "_5"%string)])]))]) |};
          {| identifier := ("merge"%string, 3) ; varl := ["_0"%string;"_1"%string;"_2"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string)]) [([(PVar "Fun"%string);(PVar "T1"%string);(PCons (PVar "H2"%string) (PVar "T2"%string))], (ETry (ELet ["_3"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_function"%string)) [(EVar "Fun"%string);(ELit (Integer (2)))]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=:="%string)) [(EVar "_3"%string);(ELit (Atom "true"%string))])) ["Try"%string] (EVar "Try"%string) ["T"%string;"R"%string] (ELit (Atom "false"%string))), (ELet ["_4"%string] (EApp (EFunId ("fmerge2_1"%string, 5)) [(EVar "T1"%string);(EVar "H2"%string);(EVar "Fun"%string);(EVar "T2"%string);ENil]) (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "_4"%string);ENil])));([(PVar "Fun"%string);(PVar "T1"%string);PNil], (ETry (ELet ["_5"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_function"%string)) [(EVar "Fun"%string);(ELit (Integer (2)))]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=:="%string)) [(EVar "_5"%string);(ELit (Atom "true"%string))])) ["Try"%string] (EVar "Try"%string) ["T"%string;"R"%string] (ELit (Atom "false"%string))), (EVar "T1"%string));([(PVar "_8"%string);(PVar "_7"%string);(PVar "_6"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_8"%string);(EVar "_7"%string);(EVar "_6"%string)])]))]) |};
          {| identifier := ("rmerge"%string, 3) ; varl := ["_0"%string;"_1"%string;"_2"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string)]) [([(PVar "Fun"%string);(PVar "T1"%string);(PCons (PVar "H2"%string) (PVar "T2"%string))], (ETry (ELet ["_3"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_function"%string)) [(EVar "Fun"%string);(ELit (Integer (2)))]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=:="%string)) [(EVar "_3"%string);(ELit (Atom "true"%string))])) ["Try"%string] (EVar "Try"%string) ["T"%string;"R"%string] (ELit (Atom "false"%string))), (ELet ["_4"%string] (EApp (EFunId ("rfmerge2_1"%string, 5)) [(EVar "T1"%string);(EVar "H2"%string);(EVar "Fun"%string);(EVar "T2"%string);ENil]) (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "_4"%string);ENil])));([(PVar "Fun"%string);(PVar "T1"%string);PNil], (ETry (ELet ["_5"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_function"%string)) [(EVar "Fun"%string);(ELit (Integer (2)))]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=:="%string)) [(EVar "_5"%string);(ELit (Atom "true"%string))])) ["Try"%string] (EVar "Try"%string) ["T"%string;"R"%string] (ELit (Atom "false"%string))), (EVar "T1"%string));([(PVar "_8"%string);(PVar "_7"%string);(PVar "_6"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_8"%string);(EVar "_7"%string);(EVar "_6"%string)])]))]) |};
          {| identifier := ("usort"%string, 2) ; varl := ["_0"%string;"_1"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string)]) [([(PVar "Fun"%string);(PTuple [(PLit (Atom "c_alias"%string));PNil;(PVar "L"%string);(PCons (PVar "_7"%string) PNil)])], (ETry (ELet ["_2"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_function"%string)) [(EVar "Fun"%string);(ELit (Integer (2)))]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=:="%string)) [(EVar "_2"%string);(ELit (Atom "true"%string))])) ["Try"%string] (EVar "Try"%string) ["T"%string;"R"%string] (ELit (Atom "false"%string))), (EVar "L"%string));([(PVar "Fun"%string);(PTuple [(PLit (Atom "c_alias"%string));PNil;(PVar "L"%string);PNil])], (ETry (ELet ["_3"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_function"%string)) [(EVar "Fun"%string);(ELit (Integer (2)))]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=:="%string)) [(EVar "_3"%string);(ELit (Atom "true"%string))])) ["Try"%string] (EVar "Try"%string) ["T"%string;"R"%string] (ELit (Atom "false"%string))), (EVar "L"%string));([(PVar "Fun"%string);(PCons (PVar "X"%string) (PVar "L"%string))], (ETry (ELet ["_4"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_function"%string)) [(EVar "Fun"%string);(ELit (Integer (2)))]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=:="%string)) [(EVar "_4"%string);(ELit (Atom "true"%string))])) ["Try"%string] (EVar "Try"%string) ["T"%string;"R"%string] (ELit (Atom "false"%string))), (EApp (EFunId ("usort_1"%string, 3)) [(EVar "Fun"%string);(EVar "X"%string);(EVar "L"%string)]));([(PVar "_6"%string);(PVar "_5"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_6"%string);(EVar "_5"%string)])]))]) |};
          {| identifier := ("usort_1"%string, 3) ; varl := ["_0"%string;"_1"%string;"_2"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string)]) [([(PVar "Fun"%string);(PVar "X"%string);(PCons (PVar "Y"%string) (PVar "L"%string))], (ELit (Atom "true"%string)), (ECase (EApp (EVar "Fun"%string) [(EVar "X"%string);(EVar "Y"%string)]) [([(PLit (Atom "true"%string))], (ELit (Atom "true"%string)), (ECase (EApp (EVar "Fun"%string) [(EVar "Y"%string);(EVar "X"%string)]) [([(PLit (Atom "true"%string))], (ELit (Atom "true"%string)), (ECase (EVar "L"%string) [([PNil], (ELit (Atom "true"%string)), (ECons (EVar "X"%string) ENil));([(PVar "_9"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("usort_1"%string, 3)) [(EVar "Fun"%string);(EVar "X"%string);(EVar "L"%string)]))]));([(PLit (Atom "false"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("ufsplit_1"%string, 6)) [(EVar "Y"%string);(EVar "X"%string);(EVar "Fun"%string);(EVar "L"%string);ENil;ENil]));([(PVar "_4"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "case_clause"%string));(EVar "_4"%string)])]))]));([(PLit (Atom "false"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("ufsplit_2"%string, 4)) [(EVar "Y"%string);(EVar "L"%string);(EVar "Fun"%string);(ECons (EVar "X"%string) ENil)]));([(PVar "_5"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "case_clause"%string));(EVar "_5"%string)])]))]));([(PVar "_8"%string);(PVar "_7"%string);(PVar "_6"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_8"%string);(EVar "_7"%string);(EVar "_6"%string)])]))]) |};
          {| identifier := ("umerge"%string, 3) ; varl := ["_0"%string;"_1"%string;"_2"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string)]) [([(PVar "Fun"%string);PNil;(PVar "T2"%string)], (ETry (ELet ["_3"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_function"%string)) [(EVar "Fun"%string);(ELit (Integer (2)))]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=:="%string)) [(EVar "_3"%string);(ELit (Atom "true"%string))])) ["Try"%string] (EVar "Try"%string) ["T"%string;"R"%string] (ELit (Atom "false"%string))), (EVar "T2"%string));([(PVar "Fun"%string);(PCons (PVar "H1"%string) (PVar "T1"%string));(PVar "T2"%string)], (ETry (ELet ["_4"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_function"%string)) [(EVar "Fun"%string);(ELit (Integer (2)))]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=:="%string)) [(EVar "_4"%string);(ELit (Atom "true"%string))])) ["Try"%string] (EVar "Try"%string) ["T"%string;"R"%string] (ELit (Atom "false"%string))), (ELet ["_5"%string] (EApp (EFunId ("ufmerge2_2"%string, 5)) [(EVar "H1"%string);(EVar "T1"%string);(EVar "Fun"%string);(EVar "T2"%string);ENil]) (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "_5"%string);ENil])));([(PVar "_8"%string);(PVar "_7"%string);(PVar "_6"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_8"%string);(EVar "_7"%string);(EVar "_6"%string)])]))]) |};
          {| identifier := ("rumerge"%string, 3) ; varl := ["_0"%string;"_1"%string;"_2"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string)]) [([(PVar "Fun"%string);(PVar "T1"%string);PNil], (ETry (ELet ["_3"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_function"%string)) [(EVar "Fun"%string);(ELit (Integer (2)))]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=:="%string)) [(EVar "_3"%string);(ELit (Atom "true"%string))])) ["Try"%string] (EVar "Try"%string) ["T"%string;"R"%string] (ELit (Atom "false"%string))), (EVar "T1"%string));([(PVar "Fun"%string);(PVar "T1"%string);(PCons (PVar "H2"%string) (PVar "T2"%string))], (ETry (ELet ["_4"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_function"%string)) [(EVar "Fun"%string);(ELit (Integer (2)))]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=:="%string)) [(EVar "_4"%string);(ELit (Atom "true"%string))])) ["Try"%string] (EVar "Try"%string) ["T"%string;"R"%string] (ELit (Atom "false"%string))), (ELet ["_5"%string] (EApp (EFunId ("rufmerge2_1"%string, 5)) [(EVar "T1"%string);(EVar "H2"%string);(EVar "Fun"%string);(EVar "T2"%string);ENil]) (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "_5"%string);ENil])));([(PVar "_8"%string);(PVar "_7"%string);(PVar "_6"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_8"%string);(EVar "_7"%string);(EVar "_6"%string)])]))]) |};
          {| identifier := ("usort"%string, 1) ; varl := ["_0"%string]; body := (ECase (EVar "_0"%string) [([(PTuple [(PLit (Atom "c_alias"%string));PNil;(PVar "L0"%string);(PCons (PVar "X"%string) (PCons (PVar "Y"%string) (PVar "L"%string)))])], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "<"%string)) [(EVar "X"%string);(EVar "Y"%string)]), (ECase (EVar "L"%string) [([PNil], (ELit (Atom "true"%string)), (EVar "L0"%string));([(PCons (PVar "Z"%string) PNil)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "<"%string)) [(EVar "Y"%string);(EVar "Z"%string)]), (EVar "L0"%string));([(PCons (PVar "Z"%string) PNil)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "Y"%string);(EVar "Z"%string)]), (ECons (EVar "X"%string) (ECons (EVar "Y"%string) ENil)));([(PCons (PVar "Z"%string) PNil)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "<"%string)) [(EVar "Z"%string);(EVar "X"%string)]), (ECons (EVar "Z"%string) (ECons (EVar "X"%string) (ECons (EVar "Y"%string) ENil))));([(PCons (PVar "Z"%string) PNil)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "Z"%string);(EVar "X"%string)]), (ECons (EVar "X"%string) (ECons (EVar "Y"%string) ENil)));([(PCons (PVar "Z"%string) PNil)], (ELit (Atom "true"%string)), (ECons (EVar "X"%string) (ECons (EVar "Z"%string) (ECons (EVar "Y"%string) ENil))));([(PVar "_4"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("usplit_1"%string, 5)) [(EVar "X"%string);(EVar "Y"%string);(EVar "L"%string);ENil;ENil]))]));([(PCons (PVar "X"%string) (PCons (PVar "Y"%string) (PVar "L"%string)))], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom ">"%string)) [(EVar "X"%string);(EVar "Y"%string)]), (ECase (EVar "L"%string) [([PNil], (ELit (Atom "true"%string)), (ECons (EVar "Y"%string) (ECons (EVar "X"%string) ENil)));([(PCons (PVar "Z"%string) PNil)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "<"%string)) [(EVar "X"%string);(EVar "Z"%string)]), (ECons (EVar "Y"%string) (ECons (EVar "X"%string) (EVar "L"%string))));([(PCons (PVar "Z"%string) PNil)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "X"%string);(EVar "Z"%string)]), (ECons (EVar "Y"%string) (ECons (EVar "X"%string) ENil)));([(PCons (PVar "Z"%string) PNil)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "<"%string)) [(EVar "Z"%string);(EVar "Y"%string)]), (ECons (EVar "Z"%string) (ECons (EVar "Y"%string) (ECons (EVar "X"%string) ENil))));([(PCons (PVar "Z"%string) PNil)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "Z"%string);(EVar "Y"%string)]), (ECons (EVar "Y"%string) (ECons (EVar "X"%string) ENil)));([(PCons (PVar "Z"%string) PNil)], (ELit (Atom "true"%string)), (ECons (EVar "Y"%string) (ECons (EVar "Z"%string) (ECons (EVar "X"%string) ENil))));([(PVar "_5"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("usplit_2"%string, 5)) [(EVar "X"%string);(EVar "Y"%string);(EVar "L"%string);ENil;ENil]))]));([(PCons (PVar "X"%string) (PCons (PVar "_Y"%string) (PVar "L"%string)))], (ELit (Atom "true"%string)), (EApp (EFunId ("usort_1"%string, 2)) [(EVar "X"%string);(EVar "L"%string)]));([(PTuple [(PLit (Atom "c_alias"%string));PNil;(PVar "L"%string);(PCons (PVar "_6"%string) PNil)])], (ELit (Atom "true"%string)), (EVar "L"%string));([PNil], (ELit (Atom "true"%string)), ENil);([(PVar "_3"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_3"%string)])]))]) |};
          {| identifier := ("usort_1"%string, 2) ; varl := ["_0"%string;"_1"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string)]) [([(PVar "X"%string);(PCons (PVar "Y"%string) (PVar "L"%string))], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "X"%string);(EVar "Y"%string)]), (EApp (EFunId ("usort_1"%string, 2)) [(EVar "X"%string);(EVar "L"%string)]));([(PVar "X"%string);(PCons (PVar "Y"%string) (PVar "L"%string))], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "<"%string)) [(EVar "X"%string);(EVar "Y"%string)]), (EApp (EFunId ("usplit_1"%string, 5)) [(EVar "X"%string);(EVar "Y"%string);(EVar "L"%string);ENil;ENil]));([(PVar "X"%string);(PCons (PVar "Y"%string) (PVar "L"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("usplit_2"%string, 5)) [(EVar "X"%string);(EVar "Y"%string);(EVar "L"%string);ENil;ENil]));([(PVar "X"%string);PNil], (ELit (Atom "true"%string)), (ECons (EVar "X"%string) ENil));([(PVar "_3"%string);(PVar "_2"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_3"%string);(EVar "_2"%string)])]))]) |};
          {| identifier := ("umerge"%string, 1) ; varl := ["_0"%string]; body := (EApp (EFunId ("umergel"%string, 1)) [(EVar "_0"%string)]) |};
          {| identifier := ("umerge3"%string, 3) ; varl := ["_0"%string;"_1"%string;"_2"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string)]) [([(PVar "L1"%string);PNil;(PVar "L3"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("umerge"%string, 2)) [(EVar "L1"%string);(EVar "L3"%string)]));([(PVar "L1"%string);(PVar "L2"%string);PNil], (ELit (Atom "true"%string)), (EApp (EFunId ("umerge"%string, 2)) [(EVar "L1"%string);(EVar "L2"%string)]));([(PVar "L1"%string);(PCons (PVar "H2"%string) (PVar "T2"%string));(PCons (PVar "H3"%string) (PVar "T3"%string))], (ELit (Atom "true"%string)), (ELet ["_3"%string] (EApp (EFunId ("umerge3_1"%string, 7)) [(EVar "L1"%string);(ECons (EVar "H2"%string) (EVar "H3"%string));(EVar "T2"%string);(EVar "H2"%string);ENil;(EVar "T3"%string);(EVar "H3"%string)]) (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "_3"%string);ENil])));([(PVar "_6"%string);(PVar "_5"%string);(PVar "_4"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_6"%string);(EVar "_5"%string);(EVar "_4"%string)])]))]) |};
          {| identifier := ("rumerge3"%string, 3) ; varl := ["_0"%string;"_1"%string;"_2"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string)]) [([(PVar "L1"%string);PNil;(PVar "L3"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rumerge"%string, 2)) [(EVar "L1"%string);(EVar "L3"%string)]));([(PVar "L1"%string);(PVar "L2"%string);PNil], (ELit (Atom "true"%string)), (EApp (EFunId ("rumerge"%string, 2)) [(EVar "L1"%string);(EVar "L2"%string)]));([(PVar "L1"%string);(PCons (PVar "H2"%string) (PVar "T2"%string));(PCons (PVar "H3"%string) (PVar "T3"%string))], (ELit (Atom "true"%string)), (ELet ["_3"%string] (EApp (EFunId ("rumerge3_1"%string, 6)) [(EVar "L1"%string);(EVar "T2"%string);(EVar "H2"%string);ENil;(EVar "T3"%string);(EVar "H3"%string)]) (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "_3"%string);ENil])));([(PVar "_6"%string);(PVar "_5"%string);(PVar "_4"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_6"%string);(EVar "_5"%string);(EVar "_4"%string)])]))]) |};
          {| identifier := ("umerge"%string, 2) ; varl := ["_0"%string;"_1"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string)]) [([PNil;(PVar "T2"%string)], (ELit (Atom "true"%string)), (EVar "T2"%string));([(PCons (PVar "H1"%string) (PVar "T1"%string));(PVar "T2"%string)], (ELit (Atom "true"%string)), (ELet ["_2"%string] (EApp (EFunId ("umerge2_2"%string, 4)) [(EVar "T1"%string);(EVar "T2"%string);ENil;(EVar "H1"%string)]) (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "_2"%string);ENil])));([(PVar "_4"%string);(PVar "_3"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_4"%string);(EVar "_3"%string)])]))]) |};
          {| identifier := ("rumerge"%string, 2) ; varl := ["_0"%string;"_1"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string)]) [([(PVar "T1"%string);PNil], (ELit (Atom "true"%string)), (EVar "T1"%string));([(PVar "T1"%string);(PCons (PVar "H2"%string) (PVar "T2"%string))], (ELit (Atom "true"%string)), (ELet ["_2"%string] (EApp (EFunId ("rumerge2_1"%string, 4)) [(EVar "T1"%string);(EVar "T2"%string);ENil;(EVar "H2"%string)]) (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "_2"%string);ENil])));([(PVar "_4"%string);(PVar "_3"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_4"%string);(EVar "_3"%string)])]))]) |};
          {| identifier := ("all"%string, 2) ; varl := ["_0"%string;"_1"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string)]) [([(PVar "Pred"%string);(PVar "List"%string)], (ETry (ELet ["_2"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_function"%string)) [(EVar "Pred"%string);(ELit (Integer (1)))]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=:="%string)) [(EVar "_2"%string);(ELit (Atom "true"%string))])) ["Try"%string] (EVar "Try"%string) ["T"%string;"R"%string] (ELit (Atom "false"%string))), (ECase (EVar "List"%string) [([(PCons (PVar "Hd"%string) (PVar "Tail"%string))], (ELit (Atom "true"%string)), (ECase (EApp (EVar "Pred"%string) [(EVar "Hd"%string)]) [([(PLit (Atom "true"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("all_1"%string, 2)) [(EVar "Pred"%string);(EVar "Tail"%string)]));([(PLit (Atom "false"%string))], (ELit (Atom "true"%string)), (ELit (Atom "false"%string)));([(PVar "_3"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "case_clause"%string));(EVar "_3"%string)])]))]));([PNil], (ELit (Atom "true"%string)), (ELit (Atom "true"%string)));([(PVar "_4"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "case_clause"%string));(EVar "_4"%string)])]))]));([(PVar "_6"%string);(PVar "_5"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_6"%string);(EVar "_5"%string)])]))]) |};
          {| identifier := ("all_1"%string, 2) ; varl := ["_0"%string;"_1"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string)]) [([(PVar "Pred"%string);(PCons (PVar "Hd"%string) (PVar "Tail"%string))], (ELit (Atom "true"%string)), (ECase (EApp (EVar "Pred"%string) [(EVar "Hd"%string)]) [([(PLit (Atom "true"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("all_1"%string, 2)) [(EVar "Pred"%string);(EVar "Tail"%string)]));([(PLit (Atom "false"%string))], (ELit (Atom "true"%string)), (ELit (Atom "false"%string)));([(PVar "_2"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "case_clause"%string));(EVar "_2"%string)])]))]));([(PVar "_Pred"%string);PNil], (ELit (Atom "true"%string)), (ELit (Atom "true"%string)));([(PVar "_4"%string);(PVar "_3"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_4"%string);(EVar "_3"%string)])]))]) |};
          {| identifier := ("any"%string, 2) ; varl := ["_0"%string;"_1"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string)]) [([(PVar "Pred"%string);(PVar "List"%string)], (ETry (ELet ["_2"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_function"%string)) [(EVar "Pred"%string);(ELit (Integer (1)))]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=:="%string)) [(EVar "_2"%string);(ELit (Atom "true"%string))])) ["Try"%string] (EVar "Try"%string) ["T"%string;"R"%string] (ELit (Atom "false"%string))), (ECase (EVar "List"%string) [([(PCons (PVar "Hd"%string) (PVar "Tail"%string))], (ELit (Atom "true"%string)), (ECase (EApp (EVar "Pred"%string) [(EVar "Hd"%string)]) [([(PLit (Atom "true"%string))], (ELit (Atom "true"%string)), (ELit (Atom "true"%string)));([(PLit (Atom "false"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("any_1"%string, 2)) [(EVar "Pred"%string);(EVar "Tail"%string)]));([(PVar "_3"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "case_clause"%string));(EVar "_3"%string)])]))]));([PNil], (ELit (Atom "true"%string)), (ELit (Atom "false"%string)));([(PVar "_4"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "case_clause"%string));(EVar "_4"%string)])]))]));([(PVar "_6"%string);(PVar "_5"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_6"%string);(EVar "_5"%string)])]))]) |};
          {| identifier := ("any_1"%string, 2) ; varl := ["_0"%string;"_1"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string)]) [([(PVar "Pred"%string);(PCons (PVar "Hd"%string) (PVar "Tail"%string))], (ELit (Atom "true"%string)), (ECase (EApp (EVar "Pred"%string) [(EVar "Hd"%string)]) [([(PLit (Atom "true"%string))], (ELit (Atom "true"%string)), (ELit (Atom "true"%string)));([(PLit (Atom "false"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("any_1"%string, 2)) [(EVar "Pred"%string);(EVar "Tail"%string)]));([(PVar "_2"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "case_clause"%string));(EVar "_2"%string)])]))]));([(PVar "_Pred"%string);PNil], (ELit (Atom "true"%string)), (ELit (Atom "false"%string)));([(PVar "_4"%string);(PVar "_3"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_4"%string);(EVar "_3"%string)])]))]) |};
          {| identifier := ("map"%string, 2) ; varl := ["_0"%string;"_1"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string)]) [([(PVar "F"%string);(PVar "List"%string)], (ETry (ELet ["_2"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_function"%string)) [(EVar "F"%string);(ELit (Integer (1)))]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=:="%string)) [(EVar "_2"%string);(ELit (Atom "true"%string))])) ["Try"%string] (EVar "Try"%string) ["T"%string;"R"%string] (ELit (Atom "false"%string))), (ECase (EVar "List"%string) [([(PCons (PVar "Hd"%string) (PVar "Tail"%string))], (ELit (Atom "true"%string)), (ELet ["_3"%string] (EApp (EVar "F"%string) [(EVar "Hd"%string)]) (ELet ["_4"%string] (EApp (EFunId ("map_1"%string, 2)) [(EVar "F"%string);(EVar "Tail"%string)]) (ECons (EVar "_3"%string) (EVar "_4"%string)))));([PNil], (ELit (Atom "true"%string)), ENil);([(PVar "_5"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "case_clause"%string));(EVar "_5"%string)])]))]));([(PVar "_7"%string);(PVar "_6"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_7"%string);(EVar "_6"%string)])]))]) |};
          {| identifier := ("map_1"%string, 2) ; varl := ["_0"%string;"_1"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string)]) [([(PVar "F"%string);(PCons (PVar "Hd"%string) (PVar "Tail"%string))], (ELit (Atom "true"%string)), (ELet ["_2"%string] (EApp (EVar "F"%string) [(EVar "Hd"%string)]) (ELet ["_3"%string] (EApp (EFunId ("map_1"%string, 2)) [(EVar "F"%string);(EVar "Tail"%string)]) (ECons (EVar "_2"%string) (EVar "_3"%string)))));([(PVar "_F"%string);PNil], (ELit (Atom "true"%string)), ENil);([(PVar "_5"%string);(PVar "_4"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_5"%string);(EVar "_4"%string)])]))]) |};
          {| identifier := ("flatmap"%string, 2) ; varl := ["_0"%string;"_1"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string)]) [([(PVar "F"%string);(PVar "List"%string)], (ETry (ELet ["_2"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_function"%string)) [(EVar "F"%string);(ELit (Integer (1)))]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=:="%string)) [(EVar "_2"%string);(ELit (Atom "true"%string))])) ["Try"%string] (EVar "Try"%string) ["T"%string;"R"%string] (ELit (Atom "false"%string))), (EApp (EFunId ("flatmap_1"%string, 2)) [(EVar "F"%string);(EVar "List"%string)]));([(PVar "_4"%string);(PVar "_3"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_4"%string);(EVar "_3"%string)])]))]) |};
          {| identifier := ("flatmap_1"%string, 2) ; varl := ["_0"%string;"_1"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string)]) [([(PVar "F"%string);(PCons (PVar "Hd"%string) (PVar "Tail"%string))], (ELit (Atom "true"%string)), (ELet ["_3"%string] (EApp (EVar "F"%string) [(EVar "Hd"%string)]) (ELet ["_2"%string] (EApp (EFunId ("flatmap_1"%string, 2)) [(EVar "F"%string);(EVar "Tail"%string)]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "++"%string)) [(EVar "_3"%string);(EVar "_2"%string)]))));([(PVar "_F"%string);PNil], (ELit (Atom "true"%string)), ENil);([(PVar "_5"%string);(PVar "_4"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_5"%string);(EVar "_4"%string)])]))]) |};
          {| identifier := ("foldl"%string, 3) ; varl := ["_0"%string;"_1"%string;"_2"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string)]) [([(PVar "F"%string);(PVar "Accu"%string);(PVar "List"%string)], (ETry (ELet ["_3"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_function"%string)) [(EVar "F"%string);(ELit (Integer (2)))]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=:="%string)) [(EVar "_3"%string);(ELit (Atom "true"%string))])) ["Try"%string] (EVar "Try"%string) ["T"%string;"R"%string] (ELit (Atom "false"%string))), (ECase (EVar "List"%string) [([(PCons (PVar "Hd"%string) (PVar "Tail"%string))], (ELit (Atom "true"%string)), (ELet ["_4"%string] (EApp (EVar "F"%string) [(EVar "Hd"%string);(EVar "Accu"%string)]) (EApp (EFunId ("foldl_1"%string, 3)) [(EVar "F"%string);(EVar "_4"%string);(EVar "Tail"%string)])));([PNil], (ELit (Atom "true"%string)), (EVar "Accu"%string));([(PVar "_5"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "case_clause"%string));(EVar "_5"%string)])]))]));([(PVar "_8"%string);(PVar "_7"%string);(PVar "_6"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_8"%string);(EVar "_7"%string);(EVar "_6"%string)])]))]) |};
          {| identifier := ("foldl_1"%string, 3) ; varl := ["_0"%string;"_1"%string;"_2"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string)]) [([(PVar "F"%string);(PVar "Accu"%string);(PCons (PVar "Hd"%string) (PVar "Tail"%string))], (ELit (Atom "true"%string)), (ELet ["_3"%string] (EApp (EVar "F"%string) [(EVar "Hd"%string);(EVar "Accu"%string)]) (EApp (EFunId ("foldl_1"%string, 3)) [(EVar "F"%string);(EVar "_3"%string);(EVar "Tail"%string)])));([(PVar "_F"%string);(PVar "Accu"%string);PNil], (ELit (Atom "true"%string)), (EVar "Accu"%string));([(PVar "_6"%string);(PVar "_5"%string);(PVar "_4"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_6"%string);(EVar "_5"%string);(EVar "_4"%string)])]))]) |};
          {| identifier := ("foldr"%string, 3) ; varl := ["_0"%string;"_1"%string;"_2"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string)]) [([(PVar "F"%string);(PVar "Accu"%string);(PVar "List"%string)], (ETry (ELet ["_3"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_function"%string)) [(EVar "F"%string);(ELit (Integer (2)))]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=:="%string)) [(EVar "_3"%string);(ELit (Atom "true"%string))])) ["Try"%string] (EVar "Try"%string) ["T"%string;"R"%string] (ELit (Atom "false"%string))), (EApp (EFunId ("foldr_1"%string, 3)) [(EVar "F"%string);(EVar "Accu"%string);(EVar "List"%string)]));([(PVar "_6"%string);(PVar "_5"%string);(PVar "_4"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_6"%string);(EVar "_5"%string);(EVar "_4"%string)])]))]) |};
          {| identifier := ("foldr_1"%string, 3) ; varl := ["_0"%string;"_1"%string;"_2"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string)]) [([(PVar "F"%string);(PVar "Accu"%string);(PCons (PVar "Hd"%string) (PVar "Tail"%string))], (ELit (Atom "true"%string)), (ELet ["_3"%string] (EApp (EFunId ("foldr_1"%string, 3)) [(EVar "F"%string);(EVar "Accu"%string);(EVar "Tail"%string)]) (EApp (EVar "F"%string) [(EVar "Hd"%string);(EVar "_3"%string)])));([(PVar "_F"%string);(PVar "Accu"%string);PNil], (ELit (Atom "true"%string)), (EVar "Accu"%string));([(PVar "_6"%string);(PVar "_5"%string);(PVar "_4"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_6"%string);(EVar "_5"%string);(EVar "_4"%string)])]))]) |};
          {| identifier := ("filter"%string, 2) ; varl := ["_0"%string;"_1"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string)]) [([(PVar "Pred"%string);(PVar "List"%string)], (ETry (ELet ["_2"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_function"%string)) [(EVar "Pred"%string);(ELit (Integer (1)))]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=:="%string)) [(EVar "_2"%string);(ELit (Atom "true"%string))])) ["Try"%string] (EVar "Try"%string) ["T"%string;"R"%string] (ELit (Atom "false"%string))), (ELetRec [(("lc$^0"%string, 1), (["_5"%string], (ECase (EVar "_5"%string) [([(PCons (PVar "E"%string) (PVar "_4"%string))], (ELit (Atom "true"%string)), (ECase (EApp (EVar "Pred"%string) [(EVar "E"%string)]) [([(PLit (Atom "true"%string))], (ELit (Atom "true"%string)), (ELet ["_7"%string] (EApp (EFunId ("lc$^0"%string, 1)) [(EVar "_4"%string)]) (ECons (EVar "E"%string) (EVar "_7"%string))));([(PLit (Atom "false"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("lc$^0"%string, 1)) [(EVar "_4"%string)]));([(PVar "_8"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "bad_filter"%string));(EVar "_8"%string)])]))]));([(PCons (PVar "E"%string) (PVar "_4"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("lc$^0"%string, 1)) [(EVar "_4"%string)]));([PNil], (ELit (Atom "true"%string)), ENil);([(PVar "_6"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "bad_generator"%string));(EVar "_6"%string)])]))])))] (EApp (EFunId ("lc$^0"%string, 1)) [(EVar "List"%string)])));([(PVar "_10"%string);(PVar "_9"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_10"%string);(EVar "_9"%string)])]))]) |};
          {| identifier := ("partition"%string, 2) ; varl := ["_0"%string;"_1"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string)]) [([(PVar "Pred"%string);(PVar "L"%string)], (ETry (ELet ["_2"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_function"%string)) [(EVar "Pred"%string);(ELit (Integer (1)))]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=:="%string)) [(EVar "_2"%string);(ELit (Atom "true"%string))])) ["Try"%string] (EVar "Try"%string) ["T"%string;"R"%string] (ELit (Atom "false"%string))), (EApp (EFunId ("partition_1"%string, 4)) [(EVar "Pred"%string);(EVar "L"%string);ENil;ENil]));([(PVar "_4"%string);(PVar "_3"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_4"%string);(EVar "_3"%string)])]))]) |};
          {| identifier := ("partition_1"%string, 4) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string)]) [([(PVar "Pred"%string);(PCons (PVar "H"%string) (PVar "T"%string));(PVar "As"%string);(PVar "Bs"%string)], (ELit (Atom "true"%string)), (ECase (EApp (EVar "Pred"%string) [(EVar "H"%string)]) [([(PLit (Atom "true"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("partition_1"%string, 4)) [(EVar "Pred"%string);(EVar "T"%string);(ECons (EVar "H"%string) (EVar "As"%string));(EVar "Bs"%string)]));([(PLit (Atom "false"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("partition_1"%string, 4)) [(EVar "Pred"%string);(EVar "T"%string);(EVar "As"%string);(ECons (EVar "H"%string) (EVar "Bs"%string))]));([(PVar "_4"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "case_clause"%string));(EVar "_4"%string)])]))]));([(PVar "_Pred"%string);PNil;(PVar "As"%string);(PVar "Bs"%string)], (ELit (Atom "true"%string)), (ELet ["_6"%string] (EApp (EFunId ("reverse"%string, 1)) [(EVar "As"%string)]) (ELet ["_5"%string] (EApp (EFunId ("reverse"%string, 1)) [(EVar "Bs"%string)]) (ETuple [(EVar "_6"%string);(EVar "_5"%string)]))));([(PVar "_10"%string);(PVar "_9"%string);(PVar "_8"%string);(PVar "_7"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_10"%string);(EVar "_9"%string);(EVar "_8"%string);(EVar "_7"%string)])]))]) |};
          {| identifier := ("filtermap"%string, 2) ; varl := ["_0"%string;"_1"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string)]) [([(PVar "F"%string);(PVar "List"%string)], (ETry (ELet ["_2"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_function"%string)) [(EVar "F"%string);(ELit (Integer (1)))]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=:="%string)) [(EVar "_2"%string);(ELit (Atom "true"%string))])) ["Try"%string] (EVar "Try"%string) ["T"%string;"R"%string] (ELit (Atom "false"%string))), (EApp (EFunId ("filtermap_1"%string, 2)) [(EVar "F"%string);(EVar "List"%string)]));([(PVar "_4"%string);(PVar "_3"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_4"%string);(EVar "_3"%string)])]))]) |};
          {| identifier := ("filtermap_1"%string, 2) ; varl := ["_0"%string;"_1"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string)]) [([(PVar "F"%string);(PCons (PVar "Hd"%string) (PVar "Tail"%string))], (ELit (Atom "true"%string)), (ECase (EApp (EVar "F"%string) [(EVar "Hd"%string)]) [([(PLit (Atom "true"%string))], (ELit (Atom "true"%string)), (ELet ["_2"%string] (EApp (EFunId ("filtermap_1"%string, 2)) [(EVar "F"%string);(EVar "Tail"%string)]) (ECons (EVar "Hd"%string) (EVar "_2"%string))));([(PTuple [(PLit (Atom "true"%string));(PVar "Val"%string)])], (ELit (Atom "true"%string)), (ELet ["_3"%string] (EApp (EFunId ("filtermap_1"%string, 2)) [(EVar "F"%string);(EVar "Tail"%string)]) (ECons (EVar "Val"%string) (EVar "_3"%string))));([(PLit (Atom "false"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("filtermap_1"%string, 2)) [(EVar "F"%string);(EVar "Tail"%string)]));([(PVar "_4"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "case_clause"%string));(EVar "_4"%string)])]))]));([(PVar "_F"%string);PNil], (ELit (Atom "true"%string)), ENil);([(PVar "_6"%string);(PVar "_5"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_6"%string);(EVar "_5"%string)])]))]) |};
          {| identifier := ("zf"%string, 2) ; varl := ["_0"%string;"_1"%string]; body := (EApp (EFunId ("filtermap"%string, 2)) [(EVar "_0"%string);(EVar "_1"%string)]) |};
          {| identifier := ("foreach"%string, 2) ; varl := ["_0"%string;"_1"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string)]) [([(PVar "F"%string);(PVar "List"%string)], (ETry (ELet ["_2"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_function"%string)) [(EVar "F"%string);(ELit (Integer (1)))]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=:="%string)) [(EVar "_2"%string);(ELit (Atom "true"%string))])) ["Try"%string] (EVar "Try"%string) ["T"%string;"R"%string] (ELit (Atom "false"%string))), (EApp (EFunId ("foreach_1"%string, 2)) [(EVar "F"%string);(EVar "List"%string)]));([(PVar "_4"%string);(PVar "_3"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_4"%string);(EVar "_3"%string)])]))]) |};
          {| identifier := ("foreach_1"%string, 2) ; varl := ["_0"%string;"_1"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string)]) [([(PVar "F"%string);(PCons (PVar "Hd"%string) (PVar "Tail"%string))], (ELit (Atom "true"%string)), (ESeq (EApp (EVar "F"%string) [(EVar "Hd"%string)]) (EApp (EFunId ("foreach_1"%string, 2)) [(EVar "F"%string);(EVar "Tail"%string)])));([(PVar "_F"%string);PNil], (ELit (Atom "true"%string)), (ELit (Atom "ok"%string)));([(PVar "_3"%string);(PVar "_2"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_3"%string);(EVar "_2"%string)])]))]) |};
          {| identifier := ("mapfoldl"%string, 3) ; varl := ["_0"%string;"_1"%string;"_2"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string)]) [([(PVar "F"%string);(PVar "Accu"%string);(PVar "List"%string)], (ETry (ELet ["_3"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_function"%string)) [(EVar "F"%string);(ELit (Integer (2)))]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=:="%string)) [(EVar "_3"%string);(ELit (Atom "true"%string))])) ["Try"%string] (EVar "Try"%string) ["T"%string;"R"%string] (ELit (Atom "false"%string))), (EApp (EFunId ("mapfoldl_1"%string, 3)) [(EVar "F"%string);(EVar "Accu"%string);(EVar "List"%string)]));([(PVar "_6"%string);(PVar "_5"%string);(PVar "_4"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_6"%string);(EVar "_5"%string);(EVar "_4"%string)])]))]) |};
          {| identifier := ("mapfoldl_1"%string, 3) ; varl := ["_0"%string;"_1"%string;"_2"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string)]) [([(PVar "F"%string);(PVar "Accu0"%string);(PCons (PVar "Hd"%string) (PVar "Tail"%string))], (ELit (Atom "true"%string)), (ECase (EApp (EVar "F"%string) [(EVar "Hd"%string);(EVar "Accu0"%string)]) [([(PTuple [(PVar "R"%string);(PVar "Accu1"%string)])], (ELit (Atom "true"%string)), (ECase (EApp (EFunId ("mapfoldl_1"%string, 3)) [(EVar "F"%string);(EVar "Accu1"%string);(EVar "Tail"%string)]) [([(PTuple [(PVar "Rs"%string);(PVar "Accu2"%string)])], (ELit (Atom "true"%string)), (ETuple [(ECons (EVar "R"%string) (EVar "Rs"%string));(EVar "Accu2"%string)]));([(PVar "_4"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "badmatch"%string));(EVar "_4"%string)])]))]));([(PVar "_3"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "badmatch"%string));(EVar "_3"%string)])]))]));([(PVar "_F"%string);(PVar "Accu"%string);PNil], (ELit (Atom "true"%string)), (ETuple [ENil;(EVar "Accu"%string)]));([(PVar "_7"%string);(PVar "_6"%string);(PVar "_5"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_7"%string);(EVar "_6"%string);(EVar "_5"%string)])]))]) |};
          {| identifier := ("mapfoldr"%string, 3) ; varl := ["_0"%string;"_1"%string;"_2"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string)]) [([(PVar "F"%string);(PVar "Accu"%string);(PVar "List"%string)], (ETry (ELet ["_3"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_function"%string)) [(EVar "F"%string);(ELit (Integer (2)))]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=:="%string)) [(EVar "_3"%string);(ELit (Atom "true"%string))])) ["Try"%string] (EVar "Try"%string) ["T"%string;"R"%string] (ELit (Atom "false"%string))), (EApp (EFunId ("mapfoldr_1"%string, 3)) [(EVar "F"%string);(EVar "Accu"%string);(EVar "List"%string)]));([(PVar "_6"%string);(PVar "_5"%string);(PVar "_4"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_6"%string);(EVar "_5"%string);(EVar "_4"%string)])]))]) |};
          {| identifier := ("mapfoldr_1"%string, 3) ; varl := ["_0"%string;"_1"%string;"_2"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string)]) [([(PVar "F"%string);(PVar "Accu0"%string);(PCons (PVar "Hd"%string) (PVar "Tail"%string))], (ELit (Atom "true"%string)), (ECase (EApp (EFunId ("mapfoldr_1"%string, 3)) [(EVar "F"%string);(EVar "Accu0"%string);(EVar "Tail"%string)]) [([(PTuple [(PVar "Rs"%string);(PVar "Accu1"%string)])], (ELit (Atom "true"%string)), (ECase (EApp (EVar "F"%string) [(EVar "Hd"%string);(EVar "Accu1"%string)]) [([(PTuple [(PVar "R"%string);(PVar "Accu2"%string)])], (ELit (Atom "true"%string)), (ETuple [(ECons (EVar "R"%string) (EVar "Rs"%string));(EVar "Accu2"%string)]));([(PVar "_4"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "badmatch"%string));(EVar "_4"%string)])]))]));([(PVar "_3"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "badmatch"%string));(EVar "_3"%string)])]))]));([(PVar "_F"%string);(PVar "Accu"%string);PNil], (ELit (Atom "true"%string)), (ETuple [ENil;(EVar "Accu"%string)]));([(PVar "_7"%string);(PVar "_6"%string);(PVar "_5"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_7"%string);(EVar "_6"%string);(EVar "_5"%string)])]))]) |};
          {| identifier := ("takewhile"%string, 2) ; varl := ["_0"%string;"_1"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string)]) [([(PVar "Pred"%string);(PVar "List"%string)], (ETry (ELet ["_2"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_function"%string)) [(EVar "Pred"%string);(ELit (Integer (1)))]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=:="%string)) [(EVar "_2"%string);(ELit (Atom "true"%string))])) ["Try"%string] (EVar "Try"%string) ["T"%string;"R"%string] (ELit (Atom "false"%string))), (EApp (EFunId ("takewhile_1"%string, 2)) [(EVar "Pred"%string);(EVar "List"%string)]));([(PVar "_4"%string);(PVar "_3"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_4"%string);(EVar "_3"%string)])]))]) |};
          {| identifier := ("takewhile_1"%string, 2) ; varl := ["_0"%string;"_1"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string)]) [([(PVar "Pred"%string);(PCons (PVar "Hd"%string) (PVar "Tail"%string))], (ELit (Atom "true"%string)), (ECase (EApp (EVar "Pred"%string) [(EVar "Hd"%string)]) [([(PLit (Atom "true"%string))], (ELit (Atom "true"%string)), (ELet ["_2"%string] (EApp (EFunId ("takewhile_1"%string, 2)) [(EVar "Pred"%string);(EVar "Tail"%string)]) (ECons (EVar "Hd"%string) (EVar "_2"%string))));([(PLit (Atom "false"%string))], (ELit (Atom "true"%string)), ENil);([(PVar "_3"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "case_clause"%string));(EVar "_3"%string)])]))]));([(PVar "_Pred"%string);PNil], (ELit (Atom "true"%string)), ENil);([(PVar "_5"%string);(PVar "_4"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_5"%string);(EVar "_4"%string)])]))]) |};
          {| identifier := ("dropwhile"%string, 2) ; varl := ["_0"%string;"_1"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string)]) [([(PVar "Pred"%string);(PVar "List"%string)], (ETry (ELet ["_2"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_function"%string)) [(EVar "Pred"%string);(ELit (Integer (1)))]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=:="%string)) [(EVar "_2"%string);(ELit (Atom "true"%string))])) ["Try"%string] (EVar "Try"%string) ["T"%string;"R"%string] (ELit (Atom "false"%string))), (EApp (EFunId ("dropwhile_1"%string, 2)) [(EVar "Pred"%string);(EVar "List"%string)]));([(PVar "_4"%string);(PVar "_3"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_4"%string);(EVar "_3"%string)])]))]) |};
          {| identifier := ("dropwhile_1"%string, 2) ; varl := ["_0"%string;"_1"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string)]) [([(PVar "Pred"%string);(PTuple [(PLit (Atom "c_alias"%string));PNil;(PVar "Rest"%string);(PCons (PVar "Hd"%string) (PVar "Tail"%string))])], (ELit (Atom "true"%string)), (ECase (EApp (EVar "Pred"%string) [(EVar "Hd"%string)]) [([(PLit (Atom "true"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("dropwhile_1"%string, 2)) [(EVar "Pred"%string);(EVar "Tail"%string)]));([(PLit (Atom "false"%string))], (ELit (Atom "true"%string)), (EVar "Rest"%string));([(PVar "_2"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "case_clause"%string));(EVar "_2"%string)])]))]));([(PVar "_Pred"%string);PNil], (ELit (Atom "true"%string)), ENil);([(PVar "_4"%string);(PVar "_3"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_4"%string);(EVar "_3"%string)])]))]) |};
          {| identifier := ("search"%string, 2) ; varl := ["_0"%string;"_1"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string)]) [([(PVar "Pred"%string);(PVar "List"%string)], (ETry (ELet ["_2"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_function"%string)) [(EVar "Pred"%string);(ELit (Integer (1)))]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=:="%string)) [(EVar "_2"%string);(ELit (Atom "true"%string))])) ["Try"%string] (EVar "Try"%string) ["T"%string;"R"%string] (ELit (Atom "false"%string))), (EApp (EFunId ("search_1"%string, 2)) [(EVar "Pred"%string);(EVar "List"%string)]));([(PVar "_4"%string);(PVar "_3"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_4"%string);(EVar "_3"%string)])]))]) |};
          {| identifier := ("search_1"%string, 2) ; varl := ["_0"%string;"_1"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string)]) [([(PVar "Pred"%string);(PCons (PVar "Hd"%string) (PVar "Tail"%string))], (ELit (Atom "true"%string)), (ECase (EApp (EVar "Pred"%string) [(EVar "Hd"%string)]) [([(PLit (Atom "true"%string))], (ELit (Atom "true"%string)), (ETuple [(ELit (Atom "value"%string));(EVar "Hd"%string)]));([(PLit (Atom "false"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("search_1"%string, 2)) [(EVar "Pred"%string);(EVar "Tail"%string)]));([(PVar "_2"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "case_clause"%string));(EVar "_2"%string)])]))]));([(PVar "_Pred"%string);PNil], (ELit (Atom "true"%string)), (ELit (Atom "false"%string)));([(PVar "_4"%string);(PVar "_3"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_4"%string);(EVar "_3"%string)])]))]) |};
          {| identifier := ("splitwith"%string, 2) ; varl := ["_0"%string;"_1"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string)]) [([(PVar "Pred"%string);(PVar "List"%string)], (ETry (ELet ["_2"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_function"%string)) [(EVar "Pred"%string);(ELit (Integer (1)))]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=:="%string)) [(EVar "_2"%string);(ELit (Atom "true"%string))])) ["Try"%string] (EVar "Try"%string) ["T"%string;"R"%string] (ELit (Atom "false"%string))), (EApp (EFunId ("splitwith_1"%string, 3)) [(EVar "Pred"%string);(EVar "List"%string);ENil]));([(PVar "_4"%string);(PVar "_3"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_4"%string);(EVar "_3"%string)])]))]) |};
          {| identifier := ("splitwith_1"%string, 3) ; varl := ["_0"%string;"_1"%string;"_2"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string)]) [([(PVar "Pred"%string);(PTuple [(PLit (Atom "c_alias"%string));(PCons (PTuple [(PLit (Integer (1549)));(PLit (Integer (19)))]) (PCons (PTuple [(PLit (Atom "file"%string));(PCons (PLit (Integer (47))) (PCons (PLit (Integer (85))) (PCons (PLit (Integer (115))) (PCons (PLit (Integer (101))) (PCons (PLit (Integer (114))) (PCons (PLit (Integer (115))) (PCons (PLit (Integer (47))) (PCons (PLit (Integer (103))) (PCons (PLit (Integer (121))) (PCons (PLit (Integer (117))) (PCons (PLit (Integer (114))) (PCons (PLit (Integer (105))) (PCons (PLit (Integer (47))) (PCons (PLit (Integer (68))) (PCons (PLit (Integer (111))) (PCons (PLit (Integer (99))) (PCons (PLit (Integer (117))) (PCons (PLit (Integer (109))) (PCons (PLit (Integer (101))) (PCons (PLit (Integer (110))) (PCons (PLit (Integer (116))) (PCons (PLit (Integer (115))) (PCons (PLit (Integer (47))) (PCons (PLit (Integer (111))) (PCons (PLit (Integer (115))) (PCons (PLit (Integer (107))) (PCons (PLit (Integer (111))) (PCons (PLit (Integer (108))) (PCons (PLit (Integer (97))) (PCons (PLit (Integer (47))) (PCons (PLit (Integer (72))) (PCons (PLit (Integer (65))) (PCons (PLit (Integer (82))) (PCons (PLit (Integer (80))) (PCons (PLit (Integer (47))) (PCons (PLit (Integer (111))) (PCons (PLit (Integer (116))) (PCons (PLit (Integer (112))) (PCons (PLit (Integer (45))) (PCons (PLit (Integer (109))) (PCons (PLit (Integer (97))) (PCons (PLit (Integer (115))) (PCons (PLit (Integer (116))) (PCons (PLit (Integer (101))) (PCons (PLit (Integer (114))) (PCons (PLit (Integer (47))) (PCons (PLit (Integer (108))) (PCons (PLit (Integer (105))) (PCons (PLit (Integer (98))) (PCons (PLit (Integer (47))) (PCons (PLit (Integer (115))) (PCons (PLit (Integer (116))) (PCons (PLit (Integer (100))) (PCons (PLit (Integer (108))) (PCons (PLit (Integer (105))) (PCons (PLit (Integer (98))) (PCons (PLit (Integer (47))) (PCons (PLit (Integer (115))) (PCons (PLit (Integer (114))) (PCons (PLit (Integer (99))) (PCons (PLit (Integer (47))) (PCons (PLit (Integer (108))) (PCons (PLit (Integer (105))) (PCons (PLit (Integer (115))) (PCons (PLit (Integer (116))) (PCons (PLit (Integer (115))) (PCons (PLit (Integer (46))) (PCons (PLit (Integer (101))) (PCons (PLit (Integer (114))) (PCons (PLit (Integer (108))) PNil))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))]) PNil));(PVar "@r0"%string);(PCons (PVar "Hd"%string) (PVar "Tail"%string))]);(PVar "Taken"%string)], (ELit (Atom "true"%string)), (ECase (EApp (EVar "Pred"%string) [(EVar "Hd"%string)]) [([(PLit (Atom "true"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("splitwith_1"%string, 3)) [(EVar "Pred"%string);(EVar "Tail"%string);(ECons (EVar "Hd"%string) (EVar "Taken"%string))]));([(PLit (Atom "false"%string))], (ELit (Atom "true"%string)), (ELet ["_3"%string] (EApp (EFunId ("reverse"%string, 1)) [(EVar "Taken"%string)]) (ETuple [(EVar "_3"%string);(EVar "@r0"%string)])));([(PVar "_4"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "case_clause"%string));(EVar "_4"%string)])]))]));([(PVar "_Pred"%string);PNil;(PVar "Taken"%string)], (ELit (Atom "true"%string)), (ELet ["_5"%string] (EApp (EFunId ("reverse"%string, 1)) [(EVar "Taken"%string)]) (ETuple [(EVar "_5"%string);ENil])));([(PVar "_8"%string);(PVar "_7"%string);(PVar "_6"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_8"%string);(EVar "_7"%string);(EVar "_6"%string)])]))]) |};
          {| identifier := ("split"%string, 2) ; varl := ["_0"%string;"_1"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string)]) [([(PVar "N"%string);(PVar "List"%string)], (ETry (ELet ["_2"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_integer"%string)) [(EVar "N"%string)]) (ELet ["_3"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom ">="%string)) [(EVar "N"%string);(ELit (Integer (0)))]) (ELet ["_4"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_list"%string)) [(EVar "List"%string)]) (ELet ["_5"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "and"%string)) [(EVar "_3"%string);(EVar "_4"%string)]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "and"%string)) [(EVar "_2"%string);(EVar "_5"%string)]))))) ["Try"%string] (EVar "Try"%string) ["T"%string;"R"%string] (ELit (Atom "false"%string))), (ECase (EApp (EFunId ("split"%string, 3)) [(EVar "N"%string);(EVar "List"%string);ENil]) [([(PTuple [(PLit (Atom "c_alias"%string));PNil;(PVar "Result"%string);(PTuple [(PVar "_9"%string);(PVar "_10"%string)])])], (ELit (Atom "true"%string)), (EVar "Result"%string));([(PVar "Fault"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_atom"%string)) [(EVar "Fault"%string)]), (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "error"%string)) [(EVar "Fault"%string);(ECons (EVar "N"%string) (ECons (EVar "List"%string) ENil))]));([(PVar "_6"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "case_clause"%string));(EVar "_6"%string)])]))]));([(PVar "N"%string);(PVar "List"%string)], (ELit (Atom "true"%string)), (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "error"%string)) [(ELit (Atom "badarg"%string));(ECons (EVar "N"%string) (ECons (EVar "List"%string) ENil))]))]) |};
          {| identifier := ("split"%string, 3) ; varl := ["_0"%string;"_1"%string;"_2"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string)]) [([(PLit (Integer (0)));(PVar "L"%string);(PVar "R"%string)], (ELit (Atom "true"%string)), (ELet ["_3"%string] (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "R"%string);ENil]) (ETuple [(EVar "_3"%string);(EVar "L"%string)])));([(PVar "N"%string);(PCons (PVar "H"%string) (PVar "T"%string));(PVar "R"%string)], (ELit (Atom "true"%string)), (ELet ["_4"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "-"%string)) [(EVar "N"%string);(ELit (Integer (1)))]) (EApp (EFunId ("split"%string, 3)) [(EVar "_4"%string);(EVar "T"%string);(ECons (EVar "H"%string) (EVar "R"%string))])));([(PVar "_8"%string);PNil;(PVar "_9"%string)], (ELit (Atom "true"%string)), (ELit (Atom "badarg"%string)));([(PVar "_7"%string);(PVar "_6"%string);(PVar "_5"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_7"%string);(EVar "_6"%string);(EVar "_5"%string)])]))]) |};
          {| identifier := ("join"%string, 2) ; varl := ["_0"%string;"_1"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string)]) [([(PVar "_Sep"%string);PNil], (ELit (Atom "true"%string)), ENil);([(PVar "Sep"%string);(PCons (PVar "H"%string) (PVar "T"%string))], (ELit (Atom "true"%string)), (ELet ["_2"%string] (EApp (EFunId ("join_prepend"%string, 2)) [(EVar "Sep"%string);(EVar "T"%string)]) (ECons (EVar "H"%string) (EVar "_2"%string))));([(PVar "_4"%string);(PVar "_3"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_4"%string);(EVar "_3"%string)])]))]) |};
          {| identifier := ("join_prepend"%string, 2) ; varl := ["_0"%string;"_1"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string)]) [([(PVar "_Sep"%string);PNil], (ELit (Atom "true"%string)), ENil);([(PVar "Sep"%string);(PCons (PVar "H"%string) (PVar "T"%string))], (ELit (Atom "true"%string)), (ELet ["_2"%string] (EApp (EFunId ("join_prepend"%string, 2)) [(EVar "Sep"%string);(EVar "T"%string)]) (ECons (EVar "Sep"%string) (ECons (EVar "H"%string) (EVar "_2"%string)))));([(PVar "_4"%string);(PVar "_3"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_4"%string);(EVar "_3"%string)])]))]) |};
          {| identifier := ("split_1"%string, 5) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string)]) [([(PVar "X"%string);(PVar "Y"%string);(PCons (PVar "Z"%string) (PVar "L"%string));(PVar "R"%string);(PVar "Rs"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom ">="%string)) [(EVar "Z"%string);(EVar "Y"%string)]), (EApp (EFunId ("split_1"%string, 5)) [(EVar "Y"%string);(EVar "Z"%string);(EVar "L"%string);(ECons (EVar "X"%string) (EVar "R"%string));(EVar "Rs"%string)]));([(PVar "X"%string);(PVar "Y"%string);(PCons (PVar "Z"%string) (PVar "L"%string));(PVar "R"%string);(PVar "Rs"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom ">="%string)) [(EVar "Z"%string);(EVar "X"%string)]), (EApp (EFunId ("split_1"%string, 5)) [(EVar "Z"%string);(EVar "Y"%string);(EVar "L"%string);(ECons (EVar "X"%string) (EVar "R"%string));(EVar "Rs"%string)]));([(PVar "X"%string);(PVar "Y"%string);(PCons (PVar "Z"%string) (PVar "L"%string));PNil;(PVar "Rs"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("split_1"%string, 5)) [(EVar "X"%string);(EVar "Y"%string);(EVar "L"%string);(ECons (EVar "Z"%string) ENil);(EVar "Rs"%string)]));([(PVar "X"%string);(PVar "Y"%string);(PCons (PVar "Z"%string) (PVar "L"%string));(PVar "R"%string);(PVar "Rs"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("split_1_1"%string, 6)) [(EVar "X"%string);(EVar "Y"%string);(EVar "L"%string);(EVar "R"%string);(EVar "Rs"%string);(EVar "Z"%string)]));([(PVar "X"%string);(PVar "Y"%string);PNil;(PVar "R"%string);(PVar "Rs"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rmergel"%string, 2)) [(ECons (ECons (EVar "Y"%string) (ECons (EVar "X"%string) (EVar "R"%string))) (EVar "Rs"%string));ENil]));([(PVar "_9"%string);(PVar "_8"%string);(PVar "_7"%string);(PVar "_6"%string);(PVar "_5"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_9"%string);(EVar "_8"%string);(EVar "_7"%string);(EVar "_6"%string);(EVar "_5"%string)])]))]) |};
          {| identifier := ("split_1_1"%string, 6) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string)]) [([(PVar "X"%string);(PVar "Y"%string);(PCons (PVar "Z"%string) (PVar "L"%string));(PVar "R"%string);(PVar "Rs"%string);(PVar "S"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom ">="%string)) [(EVar "Z"%string);(EVar "Y"%string)]), (EApp (EFunId ("split_1_1"%string, 6)) [(EVar "Y"%string);(EVar "Z"%string);(EVar "L"%string);(ECons (EVar "X"%string) (EVar "R"%string));(EVar "Rs"%string);(EVar "S"%string)]));([(PVar "X"%string);(PVar "Y"%string);(PCons (PVar "Z"%string) (PVar "L"%string));(PVar "R"%string);(PVar "Rs"%string);(PVar "S"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom ">="%string)) [(EVar "Z"%string);(EVar "X"%string)]), (EApp (EFunId ("split_1_1"%string, 6)) [(EVar "Z"%string);(EVar "Y"%string);(EVar "L"%string);(ECons (EVar "X"%string) (EVar "R"%string));(EVar "Rs"%string);(EVar "S"%string)]));([(PVar "X"%string);(PVar "Y"%string);(PCons (PVar "Z"%string) (PVar "L"%string));(PVar "R"%string);(PVar "Rs"%string);(PVar "S"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "S"%string);(EVar "Z"%string)]), (EApp (EFunId ("split_1"%string, 5)) [(EVar "S"%string);(EVar "Z"%string);(EVar "L"%string);ENil;(ECons (ECons (EVar "Y"%string) (ECons (EVar "X"%string) (EVar "R"%string))) (EVar "Rs"%string))]));([(PVar "X"%string);(PVar "Y"%string);(PCons (PVar "Z"%string) (PVar "L"%string));(PVar "R"%string);(PVar "Rs"%string);(PVar "S"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("split_1"%string, 5)) [(EVar "Z"%string);(EVar "S"%string);(EVar "L"%string);ENil;(ECons (ECons (EVar "Y"%string) (ECons (EVar "X"%string) (EVar "R"%string))) (EVar "Rs"%string))]));([(PVar "X"%string);(PVar "Y"%string);PNil;(PVar "R"%string);(PVar "Rs"%string);(PVar "S"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rmergel"%string, 2)) [(ECons (ECons (EVar "S"%string) ENil) (ECons (ECons (EVar "Y"%string) (ECons (EVar "X"%string) (EVar "R"%string))) (EVar "Rs"%string)));ENil]));([(PVar "_11"%string);(PVar "_10"%string);(PVar "_9"%string);(PVar "_8"%string);(PVar "_7"%string);(PVar "_6"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_11"%string);(EVar "_10"%string);(EVar "_9"%string);(EVar "_8"%string);(EVar "_7"%string);(EVar "_6"%string)])]))]) |};
          {| identifier := ("split_2"%string, 5) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string)]) [([(PVar "X"%string);(PVar "Y"%string);(PCons (PVar "Z"%string) (PVar "L"%string));(PVar "R"%string);(PVar "Rs"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "Z"%string);(EVar "Y"%string)]), (EApp (EFunId ("split_2"%string, 5)) [(EVar "Y"%string);(EVar "Z"%string);(EVar "L"%string);(ECons (EVar "X"%string) (EVar "R"%string));(EVar "Rs"%string)]));([(PVar "X"%string);(PVar "Y"%string);(PCons (PVar "Z"%string) (PVar "L"%string));(PVar "R"%string);(PVar "Rs"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "Z"%string);(EVar "X"%string)]), (EApp (EFunId ("split_2"%string, 5)) [(EVar "Z"%string);(EVar "Y"%string);(EVar "L"%string);(ECons (EVar "X"%string) (EVar "R"%string));(EVar "Rs"%string)]));([(PVar "X"%string);(PVar "Y"%string);(PCons (PVar "Z"%string) (PVar "L"%string));PNil;(PVar "Rs"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("split_2"%string, 5)) [(EVar "X"%string);(EVar "Y"%string);(EVar "L"%string);(ECons (EVar "Z"%string) ENil);(EVar "Rs"%string)]));([(PVar "X"%string);(PVar "Y"%string);(PCons (PVar "Z"%string) (PVar "L"%string));(PVar "R"%string);(PVar "Rs"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("split_2_1"%string, 6)) [(EVar "X"%string);(EVar "Y"%string);(EVar "L"%string);(EVar "R"%string);(EVar "Rs"%string);(EVar "Z"%string)]));([(PVar "X"%string);(PVar "Y"%string);PNil;(PVar "R"%string);(PVar "Rs"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("mergel"%string, 2)) [(ECons (ECons (EVar "Y"%string) (ECons (EVar "X"%string) (EVar "R"%string))) (EVar "Rs"%string));ENil]));([(PVar "_9"%string);(PVar "_8"%string);(PVar "_7"%string);(PVar "_6"%string);(PVar "_5"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_9"%string);(EVar "_8"%string);(EVar "_7"%string);(EVar "_6"%string);(EVar "_5"%string)])]))]) |};
          {| identifier := ("split_2_1"%string, 6) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string)]) [([(PVar "X"%string);(PVar "Y"%string);(PCons (PVar "Z"%string) (PVar "L"%string));(PVar "R"%string);(PVar "Rs"%string);(PVar "S"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "Z"%string);(EVar "Y"%string)]), (EApp (EFunId ("split_2_1"%string, 6)) [(EVar "Y"%string);(EVar "Z"%string);(EVar "L"%string);(ECons (EVar "X"%string) (EVar "R"%string));(EVar "Rs"%string);(EVar "S"%string)]));([(PVar "X"%string);(PVar "Y"%string);(PCons (PVar "Z"%string) (PVar "L"%string));(PVar "R"%string);(PVar "Rs"%string);(PVar "S"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "Z"%string);(EVar "X"%string)]), (EApp (EFunId ("split_2_1"%string, 6)) [(EVar "Z"%string);(EVar "Y"%string);(EVar "L"%string);(ECons (EVar "X"%string) (EVar "R"%string));(EVar "Rs"%string);(EVar "S"%string)]));([(PVar "X"%string);(PVar "Y"%string);(PCons (PVar "Z"%string) (PVar "L"%string));(PVar "R"%string);(PVar "Rs"%string);(PVar "S"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom ">"%string)) [(EVar "S"%string);(EVar "Z"%string)]), (EApp (EFunId ("split_2"%string, 5)) [(EVar "S"%string);(EVar "Z"%string);(EVar "L"%string);ENil;(ECons (ECons (EVar "Y"%string) (ECons (EVar "X"%string) (EVar "R"%string))) (EVar "Rs"%string))]));([(PVar "X"%string);(PVar "Y"%string);(PCons (PVar "Z"%string) (PVar "L"%string));(PVar "R"%string);(PVar "Rs"%string);(PVar "S"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("split_2"%string, 5)) [(EVar "Z"%string);(EVar "S"%string);(EVar "L"%string);ENil;(ECons (ECons (EVar "Y"%string) (ECons (EVar "X"%string) (EVar "R"%string))) (EVar "Rs"%string))]));([(PVar "X"%string);(PVar "Y"%string);PNil;(PVar "R"%string);(PVar "Rs"%string);(PVar "S"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("mergel"%string, 2)) [(ECons (ECons (EVar "S"%string) ENil) (ECons (ECons (EVar "Y"%string) (ECons (EVar "X"%string) (EVar "R"%string))) (EVar "Rs"%string)));ENil]));([(PVar "_11"%string);(PVar "_10"%string);(PVar "_9"%string);(PVar "_8"%string);(PVar "_7"%string);(PVar "_6"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_11"%string);(EVar "_10"%string);(EVar "_9"%string);(EVar "_8"%string);(EVar "_7"%string);(EVar "_6"%string)])]))]) |};
          {| identifier := ("mergel"%string, 2) ; varl := ["_0"%string;"_1"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string)]) [([(PCons PNil (PVar "L"%string));(PVar "Acc"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("mergel"%string, 2)) [(EVar "L"%string);(EVar "Acc"%string)]));([(PCons (PVar "T1"%string) (PCons (PCons (PVar "H2"%string) (PVar "T2"%string)) (PCons (PCons (PVar "H3"%string) (PVar "T3"%string)) (PVar "L"%string))));(PVar "Acc"%string)], (ELit (Atom "true"%string)), (ELet ["_2"%string] (EApp (EFunId ("merge3_1"%string, 6)) [(EVar "T1"%string);ENil;(EVar "H2"%string);(EVar "T2"%string);(EVar "H3"%string);(EVar "T3"%string)]) (EApp (EFunId ("mergel"%string, 2)) [(EVar "L"%string);(ECons (EVar "_2"%string) (EVar "Acc"%string))])));([(PCons (PVar "T1"%string) (PCons (PCons (PVar "H2"%string) (PVar "T2"%string)) PNil));(PVar "Acc"%string)], (ELit (Atom "true"%string)), (ELet ["_3"%string] (EApp (EFunId ("merge2_1"%string, 4)) [(EVar "T1"%string);(EVar "H2"%string);(EVar "T2"%string);ENil]) (EApp (EFunId ("rmergel"%string, 2)) [(ECons (EVar "_3"%string) (EVar "Acc"%string));ENil])));([(PCons (PVar "L"%string) PNil);PNil], (ELit (Atom "true"%string)), (EVar "L"%string));([(PCons (PVar "L"%string) PNil);(PVar "Acc"%string)], (ELit (Atom "true"%string)), (ELet ["_4"%string] (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "L"%string);ENil]) (EApp (EFunId ("rmergel"%string, 2)) [(ECons (EVar "_4"%string) (EVar "Acc"%string));ENil])));([PNil;PNil], (ELit (Atom "true"%string)), ENil);([PNil;(PVar "Acc"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rmergel"%string, 2)) [(EVar "Acc"%string);ENil]));([(PCons (PVar "A"%string) (PCons PNil (PVar "L"%string)));(PVar "Acc"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("mergel"%string, 2)) [(ECons (EVar "A"%string) (EVar "L"%string));(EVar "Acc"%string)]));([(PCons (PVar "A"%string) (PCons (PVar "B"%string) (PCons PNil (PVar "L"%string))));(PVar "Acc"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("mergel"%string, 2)) [(ECons (EVar "A"%string) (ECons (EVar "B"%string) (EVar "L"%string)));(EVar "Acc"%string)]));([(PVar "_6"%string);(PVar "_5"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_6"%string);(EVar "_5"%string)])]))]) |};
          {| identifier := ("rmergel"%string, 2) ; varl := ["_0"%string;"_1"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string)]) [([(PCons (PCons (PVar "H3"%string) (PVar "T3"%string)) (PCons (PCons (PVar "H2"%string) (PVar "T2"%string)) (PCons (PVar "T1"%string) (PVar "L"%string))));(PVar "Acc"%string)], (ELit (Atom "true"%string)), (ELet ["_2"%string] (EApp (EFunId ("rmerge3_1"%string, 6)) [(EVar "T1"%string);ENil;(EVar "H2"%string);(EVar "T2"%string);(EVar "H3"%string);(EVar "T3"%string)]) (EApp (EFunId ("rmergel"%string, 2)) [(EVar "L"%string);(ECons (EVar "_2"%string) (EVar "Acc"%string))])));([(PCons (PCons (PVar "H2"%string) (PVar "T2"%string)) (PCons (PVar "T1"%string) PNil));(PVar "Acc"%string)], (ELit (Atom "true"%string)), (ELet ["_3"%string] (EApp (EFunId ("rmerge2_1"%string, 4)) [(EVar "T1"%string);(EVar "H2"%string);(EVar "T2"%string);ENil]) (EApp (EFunId ("mergel"%string, 2)) [(ECons (EVar "_3"%string) (EVar "Acc"%string));ENil])));([(PCons (PVar "L"%string) PNil);(PVar "Acc"%string)], (ELit (Atom "true"%string)), (ELet ["_4"%string] (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "L"%string);ENil]) (EApp (EFunId ("mergel"%string, 2)) [(ECons (EVar "_4"%string) (EVar "Acc"%string));ENil])));([PNil;(PVar "Acc"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("mergel"%string, 2)) [(EVar "Acc"%string);ENil]));([(PVar "_6"%string);(PVar "_5"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_6"%string);(EVar "_5"%string)])]))]) |};
          {| identifier := ("merge3_1"%string, 6) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string)]) [([(PCons (PVar "H1"%string) (PVar "T1"%string));(PVar "M"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "H3"%string);(PVar "T3"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "H1"%string);(EVar "H2"%string)]), (ECase (EValues [(EVar "T1"%string);(EVar "H1"%string);(EVar "H2"%string);(EVar "T2"%string);(EVar "H3"%string);(EVar "T3"%string);(EVar "M"%string)]) [([(PVar "_20"%string);(PVar "_21"%string);(PVar "_22"%string);(PVar "_23"%string);(PVar "_24"%string);(PVar "_25"%string);(PVar "_26"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "_21"%string);(EVar "_24"%string)]), (EApp (EFunId ("merge3_1"%string, 6)) [(EVar "_20"%string);(ECons (EVar "_21"%string) (EVar "_26"%string));(EVar "_22"%string);(EVar "_23"%string);(EVar "_24"%string);(EVar "_25"%string)]));([(PVar "_27"%string);(PVar "_28"%string);(PVar "_29"%string);(PVar "_30"%string);(PVar "_31"%string);(PVar "_32"%string);(PVar "_33"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("merge3_12_3"%string, 6)) [(EVar "_27"%string);(EVar "_28"%string);(EVar "_29"%string);(EVar "_30"%string);(ECons (EVar "_31"%string) (EVar "_33"%string));(EVar "_32"%string)]))]));([(PCons (PVar "H1"%string) (PVar "T1"%string));(PVar "M"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "H3"%string);(PVar "T3"%string)], (ELit (Atom "true"%string)), (ECase (EValues [(EVar "T1"%string);(EVar "H1"%string);(EVar "H2"%string);(EVar "T2"%string);(EVar "H3"%string);(EVar "T3"%string);(EVar "M"%string)]) [([(PVar "_40"%string);(PVar "_41"%string);(PVar "_42"%string);(PVar "_43"%string);(PVar "_44"%string);(PVar "_45"%string);(PVar "_46"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "_42"%string);(EVar "_44"%string)]), (EApp (EFunId ("merge3_2"%string, 6)) [(EVar "_40"%string);(EVar "_41"%string);(ECons (EVar "_42"%string) (EVar "_46"%string));(EVar "_43"%string);(EVar "_44"%string);(EVar "_45"%string)]));([(PVar "_47"%string);(PVar "_48"%string);(PVar "_49"%string);(PVar "_50"%string);(PVar "_51"%string);(PVar "_52"%string);(PVar "_53"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("merge3_21_3"%string, 6)) [(EVar "_47"%string);(EVar "_48"%string);(EVar "_49"%string);(EVar "_50"%string);(ECons (EVar "_51"%string) (EVar "_53"%string));(EVar "_52"%string)]))]));([PNil;(PVar "M"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "H3"%string);(PVar "T3"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "H2"%string);(EVar "H3"%string)]), (EApp (EFunId ("merge2_1"%string, 4)) [(EVar "T2"%string);(EVar "H3"%string);(EVar "T3"%string);(ECons (EVar "H2"%string) (EVar "M"%string))]));([PNil;(PVar "M"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "H3"%string);(PVar "T3"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("merge2_2"%string, 5)) [(EVar "T2"%string);(EVar "H3"%string);(EVar "T3"%string);(EVar "M"%string);(EVar "H2"%string)]));([(PVar "_11"%string);(PVar "_10"%string);(PVar "_9"%string);(PVar "_8"%string);(PVar "_7"%string);(PVar "_6"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_11"%string);(EVar "_10"%string);(EVar "_9"%string);(EVar "_8"%string);(EVar "_7"%string);(EVar "_6"%string)])]))]) |};
          {| identifier := ("merge3_2"%string, 6) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string)]) [([(PVar "T1"%string);(PVar "H1"%string);(PVar "M"%string);(PCons (PVar "H2"%string) (PVar "T2"%string));(PVar "H3"%string);(PVar "T3"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "H1"%string);(EVar "H2"%string)]), (ECase (EValues [(EVar "T1"%string);(EVar "H1"%string);(EVar "H2"%string);(EVar "T2"%string);(EVar "H3"%string);(EVar "T3"%string);(EVar "M"%string)]) [([(PVar "_20"%string);(PVar "_21"%string);(PVar "_22"%string);(PVar "_23"%string);(PVar "_24"%string);(PVar "_25"%string);(PVar "_26"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "_21"%string);(EVar "_24"%string)]), (EApp (EFunId ("merge3_1"%string, 6)) [(EVar "_20"%string);(ECons (EVar "_21"%string) (EVar "_26"%string));(EVar "_22"%string);(EVar "_23"%string);(EVar "_24"%string);(EVar "_25"%string)]));([(PVar "_27"%string);(PVar "_28"%string);(PVar "_29"%string);(PVar "_30"%string);(PVar "_31"%string);(PVar "_32"%string);(PVar "_33"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("merge3_12_3"%string, 6)) [(EVar "_27"%string);(EVar "_28"%string);(EVar "_29"%string);(EVar "_30"%string);(ECons (EVar "_31"%string) (EVar "_33"%string));(EVar "_32"%string)]))]));([(PVar "T1"%string);(PVar "H1"%string);(PVar "M"%string);(PCons (PVar "H2"%string) (PVar "T2"%string));(PVar "H3"%string);(PVar "T3"%string)], (ELit (Atom "true"%string)), (ECase (EValues [(EVar "T1"%string);(EVar "H1"%string);(EVar "H2"%string);(EVar "T2"%string);(EVar "H3"%string);(EVar "T3"%string);(EVar "M"%string)]) [([(PVar "_40"%string);(PVar "_41"%string);(PVar "_42"%string);(PVar "_43"%string);(PVar "_44"%string);(PVar "_45"%string);(PVar "_46"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "_42"%string);(EVar "_44"%string)]), (EApp (EFunId ("merge3_2"%string, 6)) [(EVar "_40"%string);(EVar "_41"%string);(ECons (EVar "_42"%string) (EVar "_46"%string));(EVar "_43"%string);(EVar "_44"%string);(EVar "_45"%string)]));([(PVar "_47"%string);(PVar "_48"%string);(PVar "_49"%string);(PVar "_50"%string);(PVar "_51"%string);(PVar "_52"%string);(PVar "_53"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("merge3_21_3"%string, 6)) [(EVar "_47"%string);(EVar "_48"%string);(EVar "_49"%string);(EVar "_50"%string);(ECons (EVar "_51"%string) (EVar "_53"%string));(EVar "_52"%string)]))]));([(PVar "T1"%string);(PVar "H1"%string);(PVar "M"%string);PNil;(PVar "H3"%string);(PVar "T3"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "H1"%string);(EVar "H3"%string)]), (EApp (EFunId ("merge2_1"%string, 4)) [(EVar "T1"%string);(EVar "H3"%string);(EVar "T3"%string);(ECons (EVar "H1"%string) (EVar "M"%string))]));([(PVar "T1"%string);(PVar "H1"%string);(PVar "M"%string);PNil;(PVar "H3"%string);(PVar "T3"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("merge2_2"%string, 5)) [(EVar "T1"%string);(EVar "H3"%string);(EVar "T3"%string);(EVar "M"%string);(EVar "H1"%string)]));([(PVar "_11"%string);(PVar "_10"%string);(PVar "_9"%string);(PVar "_8"%string);(PVar "_7"%string);(PVar "_6"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_11"%string);(EVar "_10"%string);(EVar "_9"%string);(EVar "_8"%string);(EVar "_7"%string);(EVar "_6"%string)])]))]) |};
          {| identifier := ("merge3_12"%string, 7) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string;"_6"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string);(EVar "_6"%string)]) [([(PVar "T1"%string);(PVar "H1"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "H3"%string);(PVar "T3"%string);(PVar "M"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "H1"%string);(EVar "H3"%string)]), (EApp (EFunId ("merge3_1"%string, 6)) [(EVar "T1"%string);(ECons (EVar "H1"%string) (EVar "M"%string));(EVar "H2"%string);(EVar "T2"%string);(EVar "H3"%string);(EVar "T3"%string)]));([(PVar "T1"%string);(PVar "H1"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "H3"%string);(PVar "T3"%string);(PVar "M"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("merge3_12_3"%string, 6)) [(EVar "T1"%string);(EVar "H1"%string);(EVar "H2"%string);(EVar "T2"%string);(ECons (EVar "H3"%string) (EVar "M"%string));(EVar "T3"%string)]))]) |};
          {| identifier := ("merge3_12_3"%string, 6) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string)]) [([(PVar "T1"%string);(PVar "H1"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "M"%string);(PCons (PVar "H3"%string) (PVar "T3"%string))], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "H1"%string);(EVar "H3"%string)]), (EApp (EFunId ("merge3_1"%string, 6)) [(EVar "T1"%string);(ECons (EVar "H1"%string) (EVar "M"%string));(EVar "H2"%string);(EVar "T2"%string);(EVar "H3"%string);(EVar "T3"%string)]));([(PVar "T1"%string);(PVar "H1"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "M"%string);(PCons (PVar "H3"%string) (PVar "T3"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("merge3_12_3"%string, 6)) [(EVar "T1"%string);(EVar "H1"%string);(EVar "H2"%string);(EVar "T2"%string);(ECons (EVar "H3"%string) (EVar "M"%string));(EVar "T3"%string)]));([(PVar "T1"%string);(PVar "H1"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "M"%string);PNil], (ELit (Atom "true"%string)), (EApp (EFunId ("merge2_1"%string, 4)) [(EVar "T1"%string);(EVar "H2"%string);(EVar "T2"%string);(ECons (EVar "H1"%string) (EVar "M"%string))]));([(PVar "_11"%string);(PVar "_10"%string);(PVar "_9"%string);(PVar "_8"%string);(PVar "_7"%string);(PVar "_6"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_11"%string);(EVar "_10"%string);(EVar "_9"%string);(EVar "_8"%string);(EVar "_7"%string);(EVar "_6"%string)])]))]) |};
          {| identifier := ("merge3_21"%string, 7) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string;"_6"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string);(EVar "_6"%string)]) [([(PVar "T1"%string);(PVar "H1"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "H3"%string);(PVar "T3"%string);(PVar "M"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "H2"%string);(EVar "H3"%string)]), (EApp (EFunId ("merge3_2"%string, 6)) [(EVar "T1"%string);(EVar "H1"%string);(ECons (EVar "H2"%string) (EVar "M"%string));(EVar "T2"%string);(EVar "H3"%string);(EVar "T3"%string)]));([(PVar "T1"%string);(PVar "H1"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "H3"%string);(PVar "T3"%string);(PVar "M"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("merge3_21_3"%string, 6)) [(EVar "T1"%string);(EVar "H1"%string);(EVar "H2"%string);(EVar "T2"%string);(ECons (EVar "H3"%string) (EVar "M"%string));(EVar "T3"%string)]))]) |};
          {| identifier := ("merge3_21_3"%string, 6) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string)]) [([(PVar "T1"%string);(PVar "H1"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "M"%string);(PCons (PVar "H3"%string) (PVar "T3"%string))], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "H2"%string);(EVar "H3"%string)]), (EApp (EFunId ("merge3_2"%string, 6)) [(EVar "T1"%string);(EVar "H1"%string);(ECons (EVar "H2"%string) (EVar "M"%string));(EVar "T2"%string);(EVar "H3"%string);(EVar "T3"%string)]));([(PVar "T1"%string);(PVar "H1"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "M"%string);(PCons (PVar "H3"%string) (PVar "T3"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("merge3_21_3"%string, 6)) [(EVar "T1"%string);(EVar "H1"%string);(EVar "H2"%string);(EVar "T2"%string);(ECons (EVar "H3"%string) (EVar "M"%string));(EVar "T3"%string)]));([(PVar "T1"%string);(PVar "H1"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "M"%string);PNil], (ELit (Atom "true"%string)), (EApp (EFunId ("merge2_2"%string, 5)) [(EVar "T1"%string);(EVar "H2"%string);(EVar "T2"%string);(EVar "M"%string);(EVar "H1"%string)]));([(PVar "_11"%string);(PVar "_10"%string);(PVar "_9"%string);(PVar "_8"%string);(PVar "_7"%string);(PVar "_6"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_11"%string);(EVar "_10"%string);(EVar "_9"%string);(EVar "_8"%string);(EVar "_7"%string);(EVar "_6"%string)])]))]) |};
          {| identifier := ("rmerge3_1"%string, 6) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string)]) [([(PCons (PVar "H1"%string) (PVar "T1"%string));(PVar "M"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "H3"%string);(PVar "T3"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "H1"%string);(EVar "H2"%string)]), (ECase (EValues [(EVar "T1"%string);(EVar "H1"%string);(EVar "H2"%string);(EVar "T2"%string);(EVar "H3"%string);(EVar "T3"%string);(EVar "M"%string)]) [([(PVar "_20"%string);(PVar "_21"%string);(PVar "_22"%string);(PVar "_23"%string);(PVar "_24"%string);(PVar "_25"%string);(PVar "_26"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "_22"%string);(EVar "_24"%string)]), (EApp (EFunId ("rmerge3_12_3"%string, 6)) [(EVar "_20"%string);(EVar "_21"%string);(EVar "_22"%string);(EVar "_23"%string);(ECons (EVar "_24"%string) (EVar "_26"%string));(EVar "_25"%string)]));([(PVar "_27"%string);(PVar "_28"%string);(PVar "_29"%string);(PVar "_30"%string);(PVar "_31"%string);(PVar "_32"%string);(PVar "_33"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rmerge3_2"%string, 6)) [(EVar "_27"%string);(EVar "_28"%string);(ECons (EVar "_29"%string) (EVar "_33"%string));(EVar "_30"%string);(EVar "_31"%string);(EVar "_32"%string)]))]));([(PCons (PVar "H1"%string) (PVar "T1"%string));(PVar "M"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "H3"%string);(PVar "T3"%string)], (ELit (Atom "true"%string)), (ECase (EValues [(EVar "T1"%string);(EVar "H1"%string);(EVar "H2"%string);(EVar "T2"%string);(EVar "H3"%string);(EVar "T3"%string);(EVar "M"%string)]) [([(PVar "_40"%string);(PVar "_41"%string);(PVar "_42"%string);(PVar "_43"%string);(PVar "_44"%string);(PVar "_45"%string);(PVar "_46"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "_41"%string);(EVar "_44"%string)]), (EApp (EFunId ("rmerge3_21_3"%string, 6)) [(EVar "_40"%string);(EVar "_41"%string);(EVar "_42"%string);(EVar "_43"%string);(ECons (EVar "_44"%string) (EVar "_46"%string));(EVar "_45"%string)]));([(PVar "_47"%string);(PVar "_48"%string);(PVar "_49"%string);(PVar "_50"%string);(PVar "_51"%string);(PVar "_52"%string);(PVar "_53"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rmerge3_1"%string, 6)) [(EVar "_47"%string);(ECons (EVar "_48"%string) (EVar "_53"%string));(EVar "_49"%string);(EVar "_50"%string);(EVar "_51"%string);(EVar "_52"%string)]))]));([PNil;(PVar "M"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "H3"%string);(PVar "T3"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "H2"%string);(EVar "H3"%string)]), (EApp (EFunId ("rmerge2_2"%string, 5)) [(EVar "T2"%string);(EVar "H3"%string);(EVar "T3"%string);(EVar "M"%string);(EVar "H2"%string)]));([PNil;(PVar "M"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "H3"%string);(PVar "T3"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rmerge2_1"%string, 4)) [(EVar "T2"%string);(EVar "H3"%string);(EVar "T3"%string);(ECons (EVar "H2"%string) (EVar "M"%string))]));([(PVar "_11"%string);(PVar "_10"%string);(PVar "_9"%string);(PVar "_8"%string);(PVar "_7"%string);(PVar "_6"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_11"%string);(EVar "_10"%string);(EVar "_9"%string);(EVar "_8"%string);(EVar "_7"%string);(EVar "_6"%string)])]))]) |};
          {| identifier := ("rmerge3_2"%string, 6) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string)]) [([(PVar "T1"%string);(PVar "H1"%string);(PVar "M"%string);(PCons (PVar "H2"%string) (PVar "T2"%string));(PVar "H3"%string);(PVar "T3"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "H1"%string);(EVar "H2"%string)]), (ECase (EValues [(EVar "T1"%string);(EVar "H1"%string);(EVar "H2"%string);(EVar "T2"%string);(EVar "H3"%string);(EVar "T3"%string);(EVar "M"%string)]) [([(PVar "_20"%string);(PVar "_21"%string);(PVar "_22"%string);(PVar "_23"%string);(PVar "_24"%string);(PVar "_25"%string);(PVar "_26"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "_22"%string);(EVar "_24"%string)]), (EApp (EFunId ("rmerge3_12_3"%string, 6)) [(EVar "_20"%string);(EVar "_21"%string);(EVar "_22"%string);(EVar "_23"%string);(ECons (EVar "_24"%string) (EVar "_26"%string));(EVar "_25"%string)]));([(PVar "_27"%string);(PVar "_28"%string);(PVar "_29"%string);(PVar "_30"%string);(PVar "_31"%string);(PVar "_32"%string);(PVar "_33"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rmerge3_2"%string, 6)) [(EVar "_27"%string);(EVar "_28"%string);(ECons (EVar "_29"%string) (EVar "_33"%string));(EVar "_30"%string);(EVar "_31"%string);(EVar "_32"%string)]))]));([(PVar "T1"%string);(PVar "H1"%string);(PVar "M"%string);(PCons (PVar "H2"%string) (PVar "T2"%string));(PVar "H3"%string);(PVar "T3"%string)], (ELit (Atom "true"%string)), (ECase (EValues [(EVar "T1"%string);(EVar "H1"%string);(EVar "H2"%string);(EVar "T2"%string);(EVar "H3"%string);(EVar "T3"%string);(EVar "M"%string)]) [([(PVar "_40"%string);(PVar "_41"%string);(PVar "_42"%string);(PVar "_43"%string);(PVar "_44"%string);(PVar "_45"%string);(PVar "_46"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "_41"%string);(EVar "_44"%string)]), (EApp (EFunId ("rmerge3_21_3"%string, 6)) [(EVar "_40"%string);(EVar "_41"%string);(EVar "_42"%string);(EVar "_43"%string);(ECons (EVar "_44"%string) (EVar "_46"%string));(EVar "_45"%string)]));([(PVar "_47"%string);(PVar "_48"%string);(PVar "_49"%string);(PVar "_50"%string);(PVar "_51"%string);(PVar "_52"%string);(PVar "_53"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rmerge3_1"%string, 6)) [(EVar "_47"%string);(ECons (EVar "_48"%string) (EVar "_53"%string));(EVar "_49"%string);(EVar "_50"%string);(EVar "_51"%string);(EVar "_52"%string)]))]));([(PVar "T1"%string);(PVar "H1"%string);(PVar "M"%string);PNil;(PVar "H3"%string);(PVar "T3"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "H1"%string);(EVar "H3"%string)]), (EApp (EFunId ("rmerge2_2"%string, 5)) [(EVar "T1"%string);(EVar "H3"%string);(EVar "T3"%string);(EVar "M"%string);(EVar "H1"%string)]));([(PVar "T1"%string);(PVar "H1"%string);(PVar "M"%string);PNil;(PVar "H3"%string);(PVar "T3"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rmerge2_1"%string, 4)) [(EVar "T1"%string);(EVar "H3"%string);(EVar "T3"%string);(ECons (EVar "H1"%string) (EVar "M"%string))]));([(PVar "_11"%string);(PVar "_10"%string);(PVar "_9"%string);(PVar "_8"%string);(PVar "_7"%string);(PVar "_6"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_11"%string);(EVar "_10"%string);(EVar "_9"%string);(EVar "_8"%string);(EVar "_7"%string);(EVar "_6"%string)])]))]) |};
          {| identifier := ("rmerge3_12"%string, 7) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string;"_6"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string);(EVar "_6"%string)]) [([(PVar "T1"%string);(PVar "H1"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "H3"%string);(PVar "T3"%string);(PVar "M"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "H2"%string);(EVar "H3"%string)]), (EApp (EFunId ("rmerge3_12_3"%string, 6)) [(EVar "T1"%string);(EVar "H1"%string);(EVar "H2"%string);(EVar "T2"%string);(ECons (EVar "H3"%string) (EVar "M"%string));(EVar "T3"%string)]));([(PVar "T1"%string);(PVar "H1"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "H3"%string);(PVar "T3"%string);(PVar "M"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rmerge3_2"%string, 6)) [(EVar "T1"%string);(EVar "H1"%string);(ECons (EVar "H2"%string) (EVar "M"%string));(EVar "T2"%string);(EVar "H3"%string);(EVar "T3"%string)]))]) |};
          {| identifier := ("rmerge3_12_3"%string, 6) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string)]) [([(PVar "T1"%string);(PVar "H1"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "M"%string);(PCons (PVar "H3"%string) (PVar "T3"%string))], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "H2"%string);(EVar "H3"%string)]), (EApp (EFunId ("rmerge3_12_3"%string, 6)) [(EVar "T1"%string);(EVar "H1"%string);(EVar "H2"%string);(EVar "T2"%string);(ECons (EVar "H3"%string) (EVar "M"%string));(EVar "T3"%string)]));([(PVar "T1"%string);(PVar "H1"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "M"%string);(PCons (PVar "H3"%string) (PVar "T3"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("rmerge3_2"%string, 6)) [(EVar "T1"%string);(EVar "H1"%string);(ECons (EVar "H2"%string) (EVar "M"%string));(EVar "T2"%string);(EVar "H3"%string);(EVar "T3"%string)]));([(PVar "T1"%string);(PVar "H1"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "M"%string);PNil], (ELit (Atom "true"%string)), (EApp (EFunId ("rmerge2_2"%string, 5)) [(EVar "T1"%string);(EVar "H2"%string);(EVar "T2"%string);(EVar "M"%string);(EVar "H1"%string)]));([(PVar "_11"%string);(PVar "_10"%string);(PVar "_9"%string);(PVar "_8"%string);(PVar "_7"%string);(PVar "_6"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_11"%string);(EVar "_10"%string);(EVar "_9"%string);(EVar "_8"%string);(EVar "_7"%string);(EVar "_6"%string)])]))]) |};
          {| identifier := ("rmerge3_21"%string, 7) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string;"_6"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string);(EVar "_6"%string)]) [([(PVar "T1"%string);(PVar "H1"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "H3"%string);(PVar "T3"%string);(PVar "M"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "H1"%string);(EVar "H3"%string)]), (EApp (EFunId ("rmerge3_21_3"%string, 6)) [(EVar "T1"%string);(EVar "H1"%string);(EVar "H2"%string);(EVar "T2"%string);(ECons (EVar "H3"%string) (EVar "M"%string));(EVar "T3"%string)]));([(PVar "T1"%string);(PVar "H1"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "H3"%string);(PVar "T3"%string);(PVar "M"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rmerge3_1"%string, 6)) [(EVar "T1"%string);(ECons (EVar "H1"%string) (EVar "M"%string));(EVar "H2"%string);(EVar "T2"%string);(EVar "H3"%string);(EVar "T3"%string)]))]) |};
          {| identifier := ("rmerge3_21_3"%string, 6) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string)]) [([(PVar "T1"%string);(PVar "H1"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "M"%string);(PCons (PVar "H3"%string) (PVar "T3"%string))], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "H1"%string);(EVar "H3"%string)]), (EApp (EFunId ("rmerge3_21_3"%string, 6)) [(EVar "T1"%string);(EVar "H1"%string);(EVar "H2"%string);(EVar "T2"%string);(ECons (EVar "H3"%string) (EVar "M"%string));(EVar "T3"%string)]));([(PVar "T1"%string);(PVar "H1"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "M"%string);(PCons (PVar "H3"%string) (PVar "T3"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("rmerge3_1"%string, 6)) [(EVar "T1"%string);(ECons (EVar "H1"%string) (EVar "M"%string));(EVar "H2"%string);(EVar "T2"%string);(EVar "H3"%string);(EVar "T3"%string)]));([(PVar "T1"%string);(PVar "H1"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "M"%string);PNil], (ELit (Atom "true"%string)), (EApp (EFunId ("rmerge2_1"%string, 4)) [(EVar "T1"%string);(EVar "H2"%string);(EVar "T2"%string);(ECons (EVar "H1"%string) (EVar "M"%string))]));([(PVar "_11"%string);(PVar "_10"%string);(PVar "_9"%string);(PVar "_8"%string);(PVar "_7"%string);(PVar "_6"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_11"%string);(EVar "_10"%string);(EVar "_9"%string);(EVar "_8"%string);(EVar "_7"%string);(EVar "_6"%string)])]))]) |};
          {| identifier := ("merge2_1"%string, 4) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string)]) [([(PCons (PVar "H1"%string) (PVar "T1"%string));(PVar "H2"%string);(PVar "T2"%string);(PVar "M"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "H1"%string);(EVar "H2"%string)]), (EApp (EFunId ("merge2_1"%string, 4)) [(EVar "T1"%string);(EVar "H2"%string);(EVar "T2"%string);(ECons (EVar "H1"%string) (EVar "M"%string))]));([(PCons (PVar "H1"%string) (PVar "T1"%string));(PVar "H2"%string);(PVar "T2"%string);(PVar "M"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("merge2_2"%string, 5)) [(EVar "T1"%string);(EVar "H2"%string);(EVar "T2"%string);(EVar "M"%string);(EVar "H1"%string)]));([PNil;(PVar "H2"%string);(PVar "T2"%string);(PVar "M"%string)], (ELit (Atom "true"%string)), (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "T2"%string);(ECons (EVar "H2"%string) (EVar "M"%string))]));([(PVar "_7"%string);(PVar "_6"%string);(PVar "_5"%string);(PVar "_4"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_7"%string);(EVar "_6"%string);(EVar "_5"%string);(EVar "_4"%string)])]))]) |};
          {| identifier := ("merge2_2"%string, 5) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string)]) [([(PVar "T1"%string);(PVar "HdM"%string);(PCons (PVar "H2"%string) (PVar "T2"%string));(PVar "M"%string);(PVar "H1"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "H1"%string);(EVar "H2"%string)]), (EApp (EFunId ("merge2_1"%string, 4)) [(EVar "T1"%string);(EVar "H2"%string);(EVar "T2"%string);(ECons (EVar "H1"%string) (ECons (EVar "HdM"%string) (EVar "M"%string)))]));([(PVar "T1"%string);(PVar "HdM"%string);(PCons (PVar "H2"%string) (PVar "T2"%string));(PVar "M"%string);(PVar "H1"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("merge2_2"%string, 5)) [(EVar "T1"%string);(EVar "H2"%string);(EVar "T2"%string);(ECons (EVar "HdM"%string) (EVar "M"%string));(EVar "H1"%string)]));([(PVar "T1"%string);(PVar "HdM"%string);PNil;(PVar "M"%string);(PVar "H1"%string)], (ELit (Atom "true"%string)), (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "T1"%string);(ECons (EVar "H1"%string) (ECons (EVar "HdM"%string) (EVar "M"%string)))]));([(PVar "_9"%string);(PVar "_8"%string);(PVar "_7"%string);(PVar "_6"%string);(PVar "_5"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_9"%string);(EVar "_8"%string);(EVar "_7"%string);(EVar "_6"%string);(EVar "_5"%string)])]))]) |};
          {| identifier := ("rmerge2_1"%string, 4) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string)]) [([(PCons (PVar "H1"%string) (PVar "T1"%string));(PVar "H2"%string);(PVar "T2"%string);(PVar "M"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "H1"%string);(EVar "H2"%string)]), (EApp (EFunId ("rmerge2_2"%string, 5)) [(EVar "T1"%string);(EVar "H2"%string);(EVar "T2"%string);(EVar "M"%string);(EVar "H1"%string)]));([(PCons (PVar "H1"%string) (PVar "T1"%string));(PVar "H2"%string);(PVar "T2"%string);(PVar "M"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rmerge2_1"%string, 4)) [(EVar "T1"%string);(EVar "H2"%string);(EVar "T2"%string);(ECons (EVar "H1"%string) (EVar "M"%string))]));([PNil;(PVar "H2"%string);(PVar "T2"%string);(PVar "M"%string)], (ELit (Atom "true"%string)), (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "T2"%string);(ECons (EVar "H2"%string) (EVar "M"%string))]));([(PVar "_7"%string);(PVar "_6"%string);(PVar "_5"%string);(PVar "_4"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_7"%string);(EVar "_6"%string);(EVar "_5"%string);(EVar "_4"%string)])]))]) |};
          {| identifier := ("rmerge2_2"%string, 5) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string)]) [([(PVar "T1"%string);(PVar "HdM"%string);(PCons (PVar "H2"%string) (PVar "T2"%string));(PVar "M"%string);(PVar "H1"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "H1"%string);(EVar "H2"%string)]), (EApp (EFunId ("rmerge2_2"%string, 5)) [(EVar "T1"%string);(EVar "H2"%string);(EVar "T2"%string);(ECons (EVar "HdM"%string) (EVar "M"%string));(EVar "H1"%string)]));([(PVar "T1"%string);(PVar "HdM"%string);(PCons (PVar "H2"%string) (PVar "T2"%string));(PVar "M"%string);(PVar "H1"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rmerge2_1"%string, 4)) [(EVar "T1"%string);(EVar "H2"%string);(EVar "T2"%string);(ECons (EVar "H1"%string) (ECons (EVar "HdM"%string) (EVar "M"%string)))]));([(PVar "T1"%string);(PVar "HdM"%string);PNil;(PVar "M"%string);(PVar "H1"%string)], (ELit (Atom "true"%string)), (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "T1"%string);(ECons (EVar "H1"%string) (ECons (EVar "HdM"%string) (EVar "M"%string)))]));([(PVar "_9"%string);(PVar "_8"%string);(PVar "_7"%string);(PVar "_6"%string);(PVar "_5"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_9"%string);(EVar "_8"%string);(EVar "_7"%string);(EVar "_6"%string);(EVar "_5"%string)])]))]) |};
          {| identifier := ("usplit_1"%string, 5) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string)]) [([(PVar "X"%string);(PVar "Y"%string);(PCons (PVar "Z"%string) (PVar "L"%string));(PVar "R"%string);(PVar "Rs"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom ">"%string)) [(EVar "Z"%string);(EVar "Y"%string)]), (EApp (EFunId ("usplit_1"%string, 5)) [(EVar "Y"%string);(EVar "Z"%string);(EVar "L"%string);(ECons (EVar "X"%string) (EVar "R"%string));(EVar "Rs"%string)]));([(PVar "X"%string);(PVar "Y"%string);(PCons (PVar "Z"%string) (PVar "L"%string));(PVar "R"%string);(PVar "Rs"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "Z"%string);(EVar "Y"%string)]), (EApp (EFunId ("usplit_1"%string, 5)) [(EVar "X"%string);(EVar "Y"%string);(EVar "L"%string);(EVar "R"%string);(EVar "Rs"%string)]));([(PVar "X"%string);(PVar "Y"%string);(PCons (PVar "Z"%string) (PVar "L"%string));(PVar "R"%string);(PVar "Rs"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom ">"%string)) [(EVar "Z"%string);(EVar "X"%string)]), (EApp (EFunId ("usplit_1"%string, 5)) [(EVar "Z"%string);(EVar "Y"%string);(EVar "L"%string);(ECons (EVar "X"%string) (EVar "R"%string));(EVar "Rs"%string)]));([(PVar "X"%string);(PVar "Y"%string);(PCons (PVar "Z"%string) (PVar "L"%string));(PVar "R"%string);(PVar "Rs"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "Z"%string);(EVar "X"%string)]), (EApp (EFunId ("usplit_1"%string, 5)) [(EVar "X"%string);(EVar "Y"%string);(EVar "L"%string);(EVar "R"%string);(EVar "Rs"%string)]));([(PVar "X"%string);(PVar "Y"%string);(PCons (PVar "Z"%string) (PVar "L"%string));PNil;(PVar "Rs"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("usplit_1"%string, 5)) [(EVar "X"%string);(EVar "Y"%string);(EVar "L"%string);(ECons (EVar "Z"%string) ENil);(EVar "Rs"%string)]));([(PVar "X"%string);(PVar "Y"%string);(PCons (PVar "Z"%string) (PVar "L"%string));(PVar "R"%string);(PVar "Rs"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("usplit_1_1"%string, 6)) [(EVar "X"%string);(EVar "Y"%string);(EVar "L"%string);(EVar "R"%string);(EVar "Rs"%string);(EVar "Z"%string)]));([(PVar "X"%string);(PVar "Y"%string);PNil;(PVar "R"%string);(PVar "Rs"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rumergel"%string, 3)) [(ECons (ECons (EVar "Y"%string) (ECons (EVar "X"%string) (EVar "R"%string))) (EVar "Rs"%string));ENil;(ELit (Atom "asc"%string))]));([(PVar "_9"%string);(PVar "_8"%string);(PVar "_7"%string);(PVar "_6"%string);(PVar "_5"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_9"%string);(EVar "_8"%string);(EVar "_7"%string);(EVar "_6"%string);(EVar "_5"%string)])]))]) |};
          {| identifier := ("usplit_1_1"%string, 6) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string)]) [([(PVar "X"%string);(PVar "Y"%string);(PCons (PVar "Z"%string) (PVar "L"%string));(PVar "R"%string);(PVar "Rs"%string);(PVar "S"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom ">"%string)) [(EVar "Z"%string);(EVar "Y"%string)]), (EApp (EFunId ("usplit_1_1"%string, 6)) [(EVar "Y"%string);(EVar "Z"%string);(EVar "L"%string);(ECons (EVar "X"%string) (EVar "R"%string));(EVar "Rs"%string);(EVar "S"%string)]));([(PVar "X"%string);(PVar "Y"%string);(PCons (PVar "Z"%string) (PVar "L"%string));(PVar "R"%string);(PVar "Rs"%string);(PVar "S"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "Z"%string);(EVar "Y"%string)]), (EApp (EFunId ("usplit_1_1"%string, 6)) [(EVar "X"%string);(EVar "Y"%string);(EVar "L"%string);(EVar "R"%string);(EVar "Rs"%string);(EVar "S"%string)]));([(PVar "X"%string);(PVar "Y"%string);(PCons (PVar "Z"%string) (PVar "L"%string));(PVar "R"%string);(PVar "Rs"%string);(PVar "S"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom ">"%string)) [(EVar "Z"%string);(EVar "X"%string)]), (EApp (EFunId ("usplit_1_1"%string, 6)) [(EVar "Z"%string);(EVar "Y"%string);(EVar "L"%string);(ECons (EVar "X"%string) (EVar "R"%string));(EVar "Rs"%string);(EVar "S"%string)]));([(PVar "X"%string);(PVar "Y"%string);(PCons (PVar "Z"%string) (PVar "L"%string));(PVar "R"%string);(PVar "Rs"%string);(PVar "S"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "Z"%string);(EVar "X"%string)]), (EApp (EFunId ("usplit_1_1"%string, 6)) [(EVar "X"%string);(EVar "Y"%string);(EVar "L"%string);(EVar "R"%string);(EVar "Rs"%string);(EVar "S"%string)]));([(PVar "X"%string);(PVar "Y"%string);(PCons (PVar "Z"%string) (PVar "L"%string));(PVar "R"%string);(PVar "Rs"%string);(PVar "S"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom ">"%string)) [(EVar "Z"%string);(EVar "S"%string)]), (EApp (EFunId ("usplit_1"%string, 5)) [(EVar "S"%string);(EVar "Z"%string);(EVar "L"%string);ENil;(ECons (ECons (EVar "Y"%string) (ECons (EVar "X"%string) (EVar "R"%string))) (EVar "Rs"%string))]));([(PVar "X"%string);(PVar "Y"%string);(PCons (PVar "Z"%string) (PVar "L"%string));(PVar "R"%string);(PVar "Rs"%string);(PVar "S"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "Z"%string);(EVar "S"%string)]), (EApp (EFunId ("usplit_1_1"%string, 6)) [(EVar "X"%string);(EVar "Y"%string);(EVar "L"%string);(EVar "R"%string);(EVar "Rs"%string);(EVar "S"%string)]));([(PVar "X"%string);(PVar "Y"%string);(PCons (PVar "Z"%string) (PVar "L"%string));(PVar "R"%string);(PVar "Rs"%string);(PVar "S"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("usplit_1"%string, 5)) [(EVar "Z"%string);(EVar "S"%string);(EVar "L"%string);ENil;(ECons (ECons (EVar "Y"%string) (ECons (EVar "X"%string) (EVar "R"%string))) (EVar "Rs"%string))]));([(PVar "X"%string);(PVar "Y"%string);PNil;(PVar "R"%string);(PVar "Rs"%string);(PVar "S"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rumergel"%string, 3)) [(ECons (ECons (EVar "S"%string) ENil) (ECons (ECons (EVar "Y"%string) (ECons (EVar "X"%string) (EVar "R"%string))) (EVar "Rs"%string)));ENil;(ELit (Atom "asc"%string))]));([(PVar "_11"%string);(PVar "_10"%string);(PVar "_9"%string);(PVar "_8"%string);(PVar "_7"%string);(PVar "_6"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_11"%string);(EVar "_10"%string);(EVar "_9"%string);(EVar "_8"%string);(EVar "_7"%string);(EVar "_6"%string)])]))]) |};
          {| identifier := ("usplit_2"%string, 5) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string)]) [([(PVar "X"%string);(PVar "Y"%string);(PCons (PVar "Z"%string) (PVar "L"%string));(PVar "R"%string);(PVar "Rs"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "<"%string)) [(EVar "Z"%string);(EVar "Y"%string)]), (EApp (EFunId ("usplit_2"%string, 5)) [(EVar "Y"%string);(EVar "Z"%string);(EVar "L"%string);(ECons (EVar "X"%string) (EVar "R"%string));(EVar "Rs"%string)]));([(PVar "X"%string);(PVar "Y"%string);(PCons (PVar "Z"%string) (PVar "L"%string));(PVar "R"%string);(PVar "Rs"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "Z"%string);(EVar "Y"%string)]), (EApp (EFunId ("usplit_2"%string, 5)) [(EVar "X"%string);(EVar "Y"%string);(EVar "L"%string);(EVar "R"%string);(EVar "Rs"%string)]));([(PVar "X"%string);(PVar "Y"%string);(PCons (PVar "Z"%string) (PVar "L"%string));(PVar "R"%string);(PVar "Rs"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "<"%string)) [(EVar "Z"%string);(EVar "X"%string)]), (EApp (EFunId ("usplit_2"%string, 5)) [(EVar "Z"%string);(EVar "Y"%string);(EVar "L"%string);(ECons (EVar "X"%string) (EVar "R"%string));(EVar "Rs"%string)]));([(PVar "X"%string);(PVar "Y"%string);(PCons (PVar "Z"%string) (PVar "L"%string));(PVar "R"%string);(PVar "Rs"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "Z"%string);(EVar "X"%string)]), (EApp (EFunId ("usplit_2"%string, 5)) [(EVar "X"%string);(EVar "Y"%string);(EVar "L"%string);(EVar "R"%string);(EVar "Rs"%string)]));([(PVar "X"%string);(PVar "Y"%string);(PCons (PVar "Z"%string) (PVar "L"%string));PNil;(PVar "Rs"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("usplit_2"%string, 5)) [(EVar "X"%string);(EVar "Y"%string);(EVar "L"%string);(ECons (EVar "Z"%string) ENil);(EVar "Rs"%string)]));([(PVar "X"%string);(PVar "Y"%string);(PCons (PVar "Z"%string) (PVar "L"%string));(PVar "R"%string);(PVar "Rs"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("usplit_2_1"%string, 6)) [(EVar "X"%string);(EVar "Y"%string);(EVar "L"%string);(EVar "R"%string);(EVar "Rs"%string);(EVar "Z"%string)]));([(PVar "X"%string);(PVar "Y"%string);PNil;(PVar "R"%string);(PVar "Rs"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("umergel"%string, 3)) [(ECons (ECons (EVar "Y"%string) (ECons (EVar "X"%string) (EVar "R"%string))) (EVar "Rs"%string));ENil;(ELit (Atom "desc"%string))]));([(PVar "_9"%string);(PVar "_8"%string);(PVar "_7"%string);(PVar "_6"%string);(PVar "_5"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_9"%string);(EVar "_8"%string);(EVar "_7"%string);(EVar "_6"%string);(EVar "_5"%string)])]))]) |};
          {| identifier := ("usplit_2_1"%string, 6) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string)]) [([(PVar "X"%string);(PVar "Y"%string);(PCons (PVar "Z"%string) (PVar "L"%string));(PVar "R"%string);(PVar "Rs"%string);(PVar "S"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "<"%string)) [(EVar "Z"%string);(EVar "Y"%string)]), (EApp (EFunId ("usplit_2_1"%string, 6)) [(EVar "Y"%string);(EVar "Z"%string);(EVar "L"%string);(ECons (EVar "X"%string) (EVar "R"%string));(EVar "Rs"%string);(EVar "S"%string)]));([(PVar "X"%string);(PVar "Y"%string);(PCons (PVar "Z"%string) (PVar "L"%string));(PVar "R"%string);(PVar "Rs"%string);(PVar "S"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "Z"%string);(EVar "Y"%string)]), (EApp (EFunId ("usplit_2_1"%string, 6)) [(EVar "X"%string);(EVar "Y"%string);(EVar "L"%string);(EVar "R"%string);(EVar "Rs"%string);(EVar "S"%string)]));([(PVar "X"%string);(PVar "Y"%string);(PCons (PVar "Z"%string) (PVar "L"%string));(PVar "R"%string);(PVar "Rs"%string);(PVar "S"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "<"%string)) [(EVar "Z"%string);(EVar "X"%string)]), (EApp (EFunId ("usplit_2_1"%string, 6)) [(EVar "Z"%string);(EVar "Y"%string);(EVar "L"%string);(ECons (EVar "X"%string) (EVar "R"%string));(EVar "Rs"%string);(EVar "S"%string)]));([(PVar "X"%string);(PVar "Y"%string);(PCons (PVar "Z"%string) (PVar "L"%string));(PVar "R"%string);(PVar "Rs"%string);(PVar "S"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "Z"%string);(EVar "X"%string)]), (EApp (EFunId ("usplit_2_1"%string, 6)) [(EVar "X"%string);(EVar "Y"%string);(EVar "L"%string);(EVar "R"%string);(EVar "Rs"%string);(EVar "S"%string)]));([(PVar "X"%string);(PVar "Y"%string);(PCons (PVar "Z"%string) (PVar "L"%string));(PVar "R"%string);(PVar "Rs"%string);(PVar "S"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "<"%string)) [(EVar "Z"%string);(EVar "S"%string)]), (EApp (EFunId ("usplit_2"%string, 5)) [(EVar "S"%string);(EVar "Z"%string);(EVar "L"%string);ENil;(ECons (ECons (EVar "Y"%string) (ECons (EVar "X"%string) (EVar "R"%string))) (EVar "Rs"%string))]));([(PVar "X"%string);(PVar "Y"%string);(PCons (PVar "Z"%string) (PVar "L"%string));(PVar "R"%string);(PVar "Rs"%string);(PVar "S"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "Z"%string);(EVar "S"%string)]), (EApp (EFunId ("usplit_2_1"%string, 6)) [(EVar "X"%string);(EVar "Y"%string);(EVar "L"%string);(EVar "R"%string);(EVar "Rs"%string);(EVar "S"%string)]));([(PVar "X"%string);(PVar "Y"%string);(PCons (PVar "Z"%string) (PVar "L"%string));(PVar "R"%string);(PVar "Rs"%string);(PVar "S"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("usplit_2"%string, 5)) [(EVar "Z"%string);(EVar "S"%string);(EVar "L"%string);ENil;(ECons (ECons (EVar "Y"%string) (ECons (EVar "X"%string) (EVar "R"%string))) (EVar "Rs"%string))]));([(PVar "X"%string);(PVar "Y"%string);PNil;(PVar "R"%string);(PVar "Rs"%string);(PVar "S"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("umergel"%string, 3)) [(ECons (ECons (EVar "S"%string) ENil) (ECons (ECons (EVar "Y"%string) (ECons (EVar "X"%string) (EVar "R"%string))) (EVar "Rs"%string)));ENil;(ELit (Atom "desc"%string))]));([(PVar "_11"%string);(PVar "_10"%string);(PVar "_9"%string);(PVar "_8"%string);(PVar "_7"%string);(PVar "_6"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_11"%string);(EVar "_10"%string);(EVar "_9"%string);(EVar "_8"%string);(EVar "_7"%string);(EVar "_6"%string)])]))]) |};
          {| identifier := ("umergel"%string, 1) ; varl := ["_0"%string]; body := (EApp (EFunId ("umergel"%string, 3)) [(EVar "_0"%string);ENil;(ELit (Atom "asc"%string))]) |};
          {| identifier := ("umergel"%string, 3) ; varl := ["_0"%string;"_1"%string;"_2"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string)]) [([(PCons PNil (PVar "L"%string));(PVar "Acc"%string);(PVar "O"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("umergel"%string, 3)) [(EVar "L"%string);(EVar "Acc"%string);(EVar "O"%string)]));([(PCons (PVar "T1"%string) (PCons (PCons (PVar "H2"%string) (PVar "T2"%string)) (PCons (PCons (PVar "H3"%string) (PVar "T3"%string)) (PVar "L"%string))));(PVar "Acc"%string);(PLit (Atom "asc"%string))], (ELit (Atom "true"%string)), (ELet ["_3"%string] (EApp (EFunId ("umerge3_1"%string, 7)) [(EVar "T1"%string);(ECons (EVar "H2"%string) (EVar "H3"%string));(EVar "T2"%string);(EVar "H2"%string);ENil;(EVar "T3"%string);(EVar "H3"%string)]) (EApp (EFunId ("umergel"%string, 3)) [(EVar "L"%string);(ECons (EVar "_3"%string) (EVar "Acc"%string));(ELit (Atom "asc"%string))])));([(PCons (PCons (PVar "H3"%string) (PVar "T3"%string)) (PCons (PCons (PVar "H2"%string) (PVar "T2"%string)) (PCons (PVar "T1"%string) (PVar "L"%string))));(PVar "Acc"%string);(PLit (Atom "desc"%string))], (ELit (Atom "true"%string)), (ELet ["_4"%string] (EApp (EFunId ("umerge3_1"%string, 7)) [(EVar "T1"%string);(ECons (EVar "H2"%string) (EVar "H3"%string));(EVar "T2"%string);(EVar "H2"%string);ENil;(EVar "T3"%string);(EVar "H3"%string)]) (EApp (EFunId ("umergel"%string, 3)) [(EVar "L"%string);(ECons (EVar "_4"%string) (EVar "Acc"%string));(ELit (Atom "desc"%string))])));([(PCons (PVar "A"%string) (PCons PNil (PVar "L"%string)));(PVar "Acc"%string);(PVar "O"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("umergel"%string, 3)) [(ECons (EVar "A"%string) (EVar "L"%string));(EVar "Acc"%string);(EVar "O"%string)]));([(PCons (PVar "A"%string) (PCons (PVar "B"%string) (PCons PNil (PVar "L"%string))));(PVar "Acc"%string);(PVar "O"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("umergel"%string, 3)) [(ECons (EVar "A"%string) (ECons (EVar "B"%string) (EVar "L"%string)));(EVar "Acc"%string);(EVar "O"%string)]));([(PCons (PCons (PVar "H1"%string) (PVar "T1"%string)) (PCons (PVar "T2"%string) (PVar "L"%string)));(PVar "Acc"%string);(PLit (Atom "asc"%string))], (ELit (Atom "true"%string)), (ELet ["_5"%string] (EApp (EFunId ("umerge2_2"%string, 4)) [(EVar "T1"%string);(EVar "T2"%string);ENil;(EVar "H1"%string)]) (EApp (EFunId ("umergel"%string, 3)) [(EVar "L"%string);(ECons (EVar "_5"%string) (EVar "Acc"%string));(ELit (Atom "asc"%string))])));([(PCons (PVar "T2"%string) (PCons (PCons (PVar "H1"%string) (PVar "T1"%string)) (PVar "L"%string)));(PVar "Acc"%string);(PLit (Atom "desc"%string))], (ELit (Atom "true"%string)), (ELet ["_6"%string] (EApp (EFunId ("umerge2_2"%string, 4)) [(EVar "T1"%string);(EVar "T2"%string);ENil;(EVar "H1"%string)]) (EApp (EFunId ("umergel"%string, 3)) [(EVar "L"%string);(ECons (EVar "_6"%string) (EVar "Acc"%string));(ELit (Atom "desc"%string))])));([(PCons (PVar "L"%string) PNil);PNil;(PVar "_O"%string)], (ELit (Atom "true"%string)), (EVar "L"%string));([(PCons (PVar "L"%string) PNil);(PVar "Acc"%string);(PVar "O"%string)], (ELit (Atom "true"%string)), (ELet ["_7"%string] (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "L"%string);ENil]) (EApp (EFunId ("rumergel"%string, 3)) [(ECons (EVar "_7"%string) (EVar "Acc"%string));ENil;(EVar "O"%string)])));([PNil;PNil;(PVar "_O"%string)], (ELit (Atom "true"%string)), ENil);([PNil;(PVar "Acc"%string);(PVar "O"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rumergel"%string, 3)) [(EVar "Acc"%string);ENil;(EVar "O"%string)]));([(PVar "_10"%string);(PVar "_9"%string);(PVar "_8"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_10"%string);(EVar "_9"%string);(EVar "_8"%string)])]))]) |};
          {| identifier := ("rumergel"%string, 3) ; varl := ["_0"%string;"_1"%string;"_2"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string)]) [([(PCons (PCons (PVar "H3"%string) (PVar "T3"%string)) (PCons (PCons (PVar "H2"%string) (PVar "T2"%string)) (PCons (PVar "T1"%string) (PVar "L"%string))));(PVar "Acc"%string);(PLit (Atom "asc"%string))], (ELit (Atom "true"%string)), (ELet ["_3"%string] (EApp (EFunId ("rumerge3_1"%string, 6)) [(EVar "T1"%string);(EVar "T2"%string);(EVar "H2"%string);ENil;(EVar "T3"%string);(EVar "H3"%string)]) (EApp (EFunId ("rumergel"%string, 3)) [(EVar "L"%string);(ECons (EVar "_3"%string) (EVar "Acc"%string));(ELit (Atom "asc"%string))])));([(PCons (PVar "T1"%string) (PCons (PCons (PVar "H2"%string) (PVar "T2"%string)) (PCons (PCons (PVar "H3"%string) (PVar "T3"%string)) (PVar "L"%string))));(PVar "Acc"%string);(PLit (Atom "desc"%string))], (ELit (Atom "true"%string)), (ELet ["_4"%string] (EApp (EFunId ("rumerge3_1"%string, 6)) [(EVar "T1"%string);(EVar "T2"%string);(EVar "H2"%string);ENil;(EVar "T3"%string);(EVar "H3"%string)]) (EApp (EFunId ("rumergel"%string, 3)) [(EVar "L"%string);(ECons (EVar "_4"%string) (EVar "Acc"%string));(ELit (Atom "desc"%string))])));([(PCons (PCons (PVar "H2"%string) (PVar "T2"%string)) (PCons (PVar "T1"%string) (PVar "L"%string)));(PVar "Acc"%string);(PLit (Atom "asc"%string))], (ELit (Atom "true"%string)), (ELet ["_5"%string] (EApp (EFunId ("rumerge2_1"%string, 4)) [(EVar "T1"%string);(EVar "T2"%string);ENil;(EVar "H2"%string)]) (EApp (EFunId ("rumergel"%string, 3)) [(EVar "L"%string);(ECons (EVar "_5"%string) (EVar "Acc"%string));(ELit (Atom "asc"%string))])));([(PCons (PVar "T1"%string) (PCons (PCons (PVar "H2"%string) (PVar "T2"%string)) (PVar "L"%string)));(PVar "Acc"%string);(PLit (Atom "desc"%string))], (ELit (Atom "true"%string)), (ELet ["_6"%string] (EApp (EFunId ("rumerge2_1"%string, 4)) [(EVar "T1"%string);(EVar "T2"%string);ENil;(EVar "H2"%string)]) (EApp (EFunId ("rumergel"%string, 3)) [(EVar "L"%string);(ECons (EVar "_6"%string) (EVar "Acc"%string));(ELit (Atom "desc"%string))])));([(PCons (PVar "L"%string) PNil);(PVar "Acc"%string);(PVar "O"%string)], (ELit (Atom "true"%string)), (ELet ["_7"%string] (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "L"%string);ENil]) (EApp (EFunId ("umergel"%string, 3)) [(ECons (EVar "_7"%string) (EVar "Acc"%string));ENil;(EVar "O"%string)])));([PNil;(PVar "Acc"%string);(PVar "O"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("umergel"%string, 3)) [(EVar "Acc"%string);ENil;(EVar "O"%string)]));([(PVar "_10"%string);(PVar "_9"%string);(PVar "_8"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_10"%string);(EVar "_9"%string);(EVar "_8"%string)])]))]) |};
          {| identifier := ("umerge3_1"%string, 7) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string;"_6"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string);(EVar "_6"%string)]) [([(PCons (PVar "H1"%string) (PVar "T1"%string));(PVar "HdM"%string);(PVar "T2"%string);(PVar "H2"%string);(PVar "M"%string);(PVar "T3"%string);(PVar "H3"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "H1"%string);(EVar "H2"%string)]), (ECase (EValues [(EVar "T1"%string);(EVar "H1"%string);(EVar "T2"%string);(EVar "H2"%string);(EVar "M"%string);(EVar "T3"%string);(EVar "H3"%string);(EVar "HdM"%string)]) [([(PVar "_23"%string);(PVar "_24"%string);(PVar "_25"%string);(PVar "_26"%string);(PVar "_27"%string);(PVar "_28"%string);(PVar "_29"%string);(PVar "_HdM"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "_24"%string);(EVar "_29"%string)]), (EApp (EFunId ("umerge3_1"%string, 7)) [(EVar "_23"%string);(EVar "_24"%string);(EVar "_25"%string);(EVar "_26"%string);(ECons (EVar "_24"%string) (EVar "_27"%string));(EVar "_28"%string);(EVar "_29"%string)]));([(PVar "_30"%string);(PVar "_31"%string);(PVar "_32"%string);(PVar "_33"%string);(PVar "_34"%string);(PVar "_35"%string);(PVar "_36"%string);(PVar "_37"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "_36"%string);(EVar "_37"%string)]), (EApp (EFunId ("umerge3_12_3"%string, 6)) [(EVar "_30"%string);(EVar "_31"%string);(EVar "_32"%string);(EVar "_33"%string);(EVar "_34"%string);(EVar "_35"%string)]));([(PVar "_38"%string);(PVar "_39"%string);(PVar "_40"%string);(PVar "_41"%string);(PVar "_42"%string);(PVar "_43"%string);(PVar "_44"%string);(PVar "_HdM"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("umerge3_12_3"%string, 6)) [(EVar "_38"%string);(EVar "_39"%string);(EVar "_40"%string);(EVar "_41"%string);(ECons (EVar "_44"%string) (EVar "_42"%string));(EVar "_43"%string)]))]));([(PCons (PVar "H1"%string) (PVar "T1"%string));(PVar "HdM"%string);(PVar "T2"%string);(PVar "H2"%string);(PVar "M"%string);(PVar "T3"%string);(PVar "H3"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "H2"%string);(EVar "HdM"%string)]), (EApp (EFunId ("umerge3_2"%string, 7)) [(EVar "T1"%string);(EVar "H1"%string);(EVar "T2"%string);(EVar "H2"%string);(EVar "M"%string);(EVar "T3"%string);(EVar "H3"%string)]));([(PCons (PVar "H1"%string) (PVar "T1"%string));(PVar "HdM"%string);(PVar "T2"%string);(PVar "H2"%string);(PVar "M"%string);(PVar "T3"%string);(PVar "H3"%string)], (ELit (Atom "true"%string)), (ECase (EValues [(EVar "T1"%string);(EVar "H1"%string);(EVar "T2"%string);(EVar "H2"%string);(EVar "M"%string);(EVar "T3"%string);(EVar "H3"%string);(EVar "HdM"%string)]) [([(PVar "_52"%string);(PVar "_53"%string);(PVar "_54"%string);(PVar "_55"%string);(PVar "_56"%string);(PVar "_57"%string);(PVar "_58"%string);(PVar "_HdM"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "_55"%string);(EVar "_58"%string)]), (EApp (EFunId ("umerge3_2"%string, 7)) [(EVar "_52"%string);(EVar "_53"%string);(EVar "_54"%string);(EVar "_55"%string);(ECons (EVar "_55"%string) (EVar "_56"%string));(EVar "_57"%string);(EVar "_58"%string)]));([(PVar "_59"%string);(PVar "_60"%string);(PVar "_61"%string);(PVar "_62"%string);(PVar "_63"%string);(PVar "_64"%string);(PVar "_65"%string);(PVar "_66"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "_65"%string);(EVar "_66"%string)]), (EApp (EFunId ("umerge3_21_3"%string, 6)) [(EVar "_59"%string);(EVar "_60"%string);(EVar "_61"%string);(EVar "_62"%string);(EVar "_63"%string);(EVar "_64"%string)]));([(PVar "_67"%string);(PVar "_68"%string);(PVar "_69"%string);(PVar "_70"%string);(PVar "_71"%string);(PVar "_72"%string);(PVar "_73"%string);(PVar "_HdM"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("umerge3_21_3"%string, 6)) [(EVar "_67"%string);(EVar "_68"%string);(EVar "_69"%string);(EVar "_70"%string);(ECons (EVar "_73"%string) (EVar "_71"%string));(EVar "_72"%string)]))]));([PNil;(PVar "HdM"%string);(PVar "T2"%string);(PVar "H2"%string);(PVar "M"%string);(PVar "T3"%string);(PVar "H3"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "H2"%string);(EVar "HdM"%string)]), (EApp (EFunId ("umerge2_1"%string, 5)) [(EVar "T2"%string);(EVar "T3"%string);(EVar "M"%string);(EVar "HdM"%string);(EVar "H3"%string)]));([PNil;(PVar "_HdM"%string);(PVar "T2"%string);(PVar "H2"%string);(PVar "M"%string);(PVar "T3"%string);(PVar "H3"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "H2"%string);(EVar "H3"%string)]), (EApp (EFunId ("umerge2_1"%string, 5)) [(EVar "T2"%string);(EVar "T3"%string);(ECons (EVar "H2"%string) (EVar "M"%string));(EVar "H2"%string);(EVar "H3"%string)]));([PNil;(PVar "HdM"%string);(PVar "T2"%string);(PVar "H2"%string);(PVar "M"%string);(PVar "T3"%string);(PVar "H3"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "H3"%string);(EVar "HdM"%string)]), (EApp (EFunId ("umerge2_2"%string, 4)) [(EVar "T2"%string);(EVar "T3"%string);(EVar "M"%string);(EVar "H2"%string)]));([PNil;(PVar "_HdM"%string);(PVar "T2"%string);(PVar "H2"%string);(PVar "M"%string);(PVar "T3"%string);(PVar "H3"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("umerge2_2"%string, 4)) [(EVar "T2"%string);(EVar "T3"%string);(ECons (EVar "H3"%string) (EVar "M"%string));(EVar "H2"%string)]));([(PVar "_13"%string);(PVar "_12"%string);(PVar "_11"%string);(PVar "_10"%string);(PVar "_9"%string);(PVar "_8"%string);(PVar "_7"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_13"%string);(EVar "_12"%string);(EVar "_11"%string);(EVar "_10"%string);(EVar "_9"%string);(EVar "_8"%string);(EVar "_7"%string)])]))]) |};
          {| identifier := ("umerge3_2"%string, 7) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string;"_6"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string);(EVar "_6"%string)]) [([(PVar "T1"%string);(PVar "H1"%string);(PCons (PVar "H2"%string) (PVar "T2"%string));(PVar "HdM"%string);(PVar "M"%string);(PVar "T3"%string);(PVar "H3"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "H1"%string);(EVar "H2"%string)]), (ECase (EValues [(EVar "T1"%string);(EVar "H1"%string);(EVar "T2"%string);(EVar "H2"%string);(EVar "M"%string);(EVar "T3"%string);(EVar "H3"%string);(EVar "HdM"%string)]) [([(PVar "_23"%string);(PVar "_24"%string);(PVar "_25"%string);(PVar "_26"%string);(PVar "_27"%string);(PVar "_28"%string);(PVar "_29"%string);(PVar "_HdM"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "_24"%string);(EVar "_29"%string)]), (EApp (EFunId ("umerge3_1"%string, 7)) [(EVar "_23"%string);(EVar "_24"%string);(EVar "_25"%string);(EVar "_26"%string);(ECons (EVar "_24"%string) (EVar "_27"%string));(EVar "_28"%string);(EVar "_29"%string)]));([(PVar "_30"%string);(PVar "_31"%string);(PVar "_32"%string);(PVar "_33"%string);(PVar "_34"%string);(PVar "_35"%string);(PVar "_36"%string);(PVar "_37"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "_36"%string);(EVar "_37"%string)]), (EApp (EFunId ("umerge3_12_3"%string, 6)) [(EVar "_30"%string);(EVar "_31"%string);(EVar "_32"%string);(EVar "_33"%string);(EVar "_34"%string);(EVar "_35"%string)]));([(PVar "_38"%string);(PVar "_39"%string);(PVar "_40"%string);(PVar "_41"%string);(PVar "_42"%string);(PVar "_43"%string);(PVar "_44"%string);(PVar "_HdM"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("umerge3_12_3"%string, 6)) [(EVar "_38"%string);(EVar "_39"%string);(EVar "_40"%string);(EVar "_41"%string);(ECons (EVar "_44"%string) (EVar "_42"%string));(EVar "_43"%string)]))]));([(PVar "T1"%string);(PVar "H1"%string);(PCons (PVar "H2"%string) (PVar "T2"%string));(PVar "HdM"%string);(PVar "M"%string);(PVar "T3"%string);(PVar "H3"%string)], (ELit (Atom "true"%string)), (ECase (EValues [(EVar "T1"%string);(EVar "H1"%string);(EVar "T2"%string);(EVar "H2"%string);(EVar "M"%string);(EVar "T3"%string);(EVar "H3"%string);(EVar "HdM"%string)]) [([(PVar "_52"%string);(PVar "_53"%string);(PVar "_54"%string);(PVar "_55"%string);(PVar "_56"%string);(PVar "_57"%string);(PVar "_58"%string);(PVar "_HdM"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "_55"%string);(EVar "_58"%string)]), (EApp (EFunId ("umerge3_2"%string, 7)) [(EVar "_52"%string);(EVar "_53"%string);(EVar "_54"%string);(EVar "_55"%string);(ECons (EVar "_55"%string) (EVar "_56"%string));(EVar "_57"%string);(EVar "_58"%string)]));([(PVar "_59"%string);(PVar "_60"%string);(PVar "_61"%string);(PVar "_62"%string);(PVar "_63"%string);(PVar "_64"%string);(PVar "_65"%string);(PVar "_66"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "_65"%string);(EVar "_66"%string)]), (EApp (EFunId ("umerge3_21_3"%string, 6)) [(EVar "_59"%string);(EVar "_60"%string);(EVar "_61"%string);(EVar "_62"%string);(EVar "_63"%string);(EVar "_64"%string)]));([(PVar "_67"%string);(PVar "_68"%string);(PVar "_69"%string);(PVar "_70"%string);(PVar "_71"%string);(PVar "_72"%string);(PVar "_73"%string);(PVar "_HdM"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("umerge3_21_3"%string, 6)) [(EVar "_67"%string);(EVar "_68"%string);(EVar "_69"%string);(EVar "_70"%string);(ECons (EVar "_73"%string) (EVar "_71"%string));(EVar "_72"%string)]))]));([(PVar "T1"%string);(PVar "H1"%string);PNil;(PVar "_HdM"%string);(PVar "M"%string);(PVar "T3"%string);(PVar "H3"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "H1"%string);(EVar "H3"%string)]), (EApp (EFunId ("umerge2_1"%string, 5)) [(EVar "T1"%string);(EVar "T3"%string);(ECons (EVar "H1"%string) (EVar "M"%string));(EVar "H1"%string);(EVar "H3"%string)]));([(PVar "T1"%string);(PVar "H1"%string);PNil;(PVar "HdM"%string);(PVar "M"%string);(PVar "T3"%string);(PVar "H3"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "H3"%string);(EVar "HdM"%string)]), (EApp (EFunId ("umerge2_2"%string, 4)) [(EVar "T1"%string);(EVar "T3"%string);(EVar "M"%string);(EVar "H1"%string)]));([(PVar "T1"%string);(PVar "H1"%string);PNil;(PVar "_HdM"%string);(PVar "M"%string);(PVar "T3"%string);(PVar "H3"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("umerge2_2"%string, 4)) [(EVar "T1"%string);(EVar "T3"%string);(ECons (EVar "H3"%string) (EVar "M"%string));(EVar "H1"%string)]));([(PVar "_13"%string);(PVar "_12"%string);(PVar "_11"%string);(PVar "_10"%string);(PVar "_9"%string);(PVar "_8"%string);(PVar "_7"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_13"%string);(EVar "_12"%string);(EVar "_11"%string);(EVar "_10"%string);(EVar "_9"%string);(EVar "_8"%string);(EVar "_7"%string)])]))]) |};
          {| identifier := ("umerge3_12"%string, 8) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string;"_6"%string;"_7"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string);(EVar "_6"%string);(EVar "_7"%string)]) [([(PVar "T1"%string);(PVar "H1"%string);(PVar "T2"%string);(PVar "H2"%string);(PVar "M"%string);(PVar "T3"%string);(PVar "H3"%string);(PVar "_HdM"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "H1"%string);(EVar "H3"%string)]), (EApp (EFunId ("umerge3_1"%string, 7)) [(EVar "T1"%string);(EVar "H1"%string);(EVar "T2"%string);(EVar "H2"%string);(ECons (EVar "H1"%string) (EVar "M"%string));(EVar "T3"%string);(EVar "H3"%string)]));([(PVar "T1"%string);(PVar "H1"%string);(PVar "T2"%string);(PVar "H2"%string);(PVar "M"%string);(PVar "T3"%string);(PVar "H3"%string);(PVar "HdM"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "H3"%string);(EVar "HdM"%string)]), (EApp (EFunId ("umerge3_12_3"%string, 6)) [(EVar "T1"%string);(EVar "H1"%string);(EVar "T2"%string);(EVar "H2"%string);(EVar "M"%string);(EVar "T3"%string)]));([(PVar "T1"%string);(PVar "H1"%string);(PVar "T2"%string);(PVar "H2"%string);(PVar "M"%string);(PVar "T3"%string);(PVar "H3"%string);(PVar "_HdM"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("umerge3_12_3"%string, 6)) [(EVar "T1"%string);(EVar "H1"%string);(EVar "T2"%string);(EVar "H2"%string);(ECons (EVar "H3"%string) (EVar "M"%string));(EVar "T3"%string)]))]) |};
          {| identifier := ("umerge3_12_3"%string, 6) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string)]) [([(PVar "T1"%string);(PVar "H1"%string);(PVar "T2"%string);(PVar "H2"%string);(PVar "M"%string);(PCons (PVar "H3"%string) (PVar "T3"%string))], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "H1"%string);(EVar "H3"%string)]), (EApp (EFunId ("umerge3_1"%string, 7)) [(EVar "T1"%string);(EVar "H1"%string);(EVar "T2"%string);(EVar "H2"%string);(ECons (EVar "H1"%string) (EVar "M"%string));(EVar "T3"%string);(EVar "H3"%string)]));([(PVar "T1"%string);(PVar "H1"%string);(PVar "T2"%string);(PVar "H2"%string);(PVar "M"%string);(PCons (PVar "H3"%string) (PVar "T3"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("umerge3_12_3"%string, 6)) [(EVar "T1"%string);(EVar "H1"%string);(EVar "T2"%string);(EVar "H2"%string);(ECons (EVar "H3"%string) (EVar "M"%string));(EVar "T3"%string)]));([(PVar "T1"%string);(PVar "H1"%string);(PVar "T2"%string);(PVar "H2"%string);(PVar "M"%string);PNil], (ELit (Atom "true"%string)), (EApp (EFunId ("umerge2_1"%string, 5)) [(EVar "T1"%string);(EVar "T2"%string);(ECons (EVar "H1"%string) (EVar "M"%string));(EVar "H1"%string);(EVar "H2"%string)]));([(PVar "_11"%string);(PVar "_10"%string);(PVar "_9"%string);(PVar "_8"%string);(PVar "_7"%string);(PVar "_6"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_11"%string);(EVar "_10"%string);(EVar "_9"%string);(EVar "_8"%string);(EVar "_7"%string);(EVar "_6"%string)])]))]) |};
          {| identifier := ("umerge3_21"%string, 8) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string;"_6"%string;"_7"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string);(EVar "_6"%string);(EVar "_7"%string)]) [([(PVar "T1"%string);(PVar "H1"%string);(PVar "T2"%string);(PVar "H2"%string);(PVar "M"%string);(PVar "T3"%string);(PVar "H3"%string);(PVar "_HdM"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "H2"%string);(EVar "H3"%string)]), (EApp (EFunId ("umerge3_2"%string, 7)) [(EVar "T1"%string);(EVar "H1"%string);(EVar "T2"%string);(EVar "H2"%string);(ECons (EVar "H2"%string) (EVar "M"%string));(EVar "T3"%string);(EVar "H3"%string)]));([(PVar "T1"%string);(PVar "H1"%string);(PVar "T2"%string);(PVar "H2"%string);(PVar "M"%string);(PVar "T3"%string);(PVar "H3"%string);(PVar "HdM"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "H3"%string);(EVar "HdM"%string)]), (EApp (EFunId ("umerge3_21_3"%string, 6)) [(EVar "T1"%string);(EVar "H1"%string);(EVar "T2"%string);(EVar "H2"%string);(EVar "M"%string);(EVar "T3"%string)]));([(PVar "T1"%string);(PVar "H1"%string);(PVar "T2"%string);(PVar "H2"%string);(PVar "M"%string);(PVar "T3"%string);(PVar "H3"%string);(PVar "_HdM"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("umerge3_21_3"%string, 6)) [(EVar "T1"%string);(EVar "H1"%string);(EVar "T2"%string);(EVar "H2"%string);(ECons (EVar "H3"%string) (EVar "M"%string));(EVar "T3"%string)]))]) |};
          {| identifier := ("umerge3_21_3"%string, 6) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string)]) [([(PVar "T1"%string);(PVar "H1"%string);(PVar "T2"%string);(PVar "H2"%string);(PVar "M"%string);(PCons (PVar "H3"%string) (PVar "T3"%string))], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "H2"%string);(EVar "H3"%string)]), (EApp (EFunId ("umerge3_2"%string, 7)) [(EVar "T1"%string);(EVar "H1"%string);(EVar "T2"%string);(EVar "H2"%string);(ECons (EVar "H2"%string) (EVar "M"%string));(EVar "T3"%string);(EVar "H3"%string)]));([(PVar "T1"%string);(PVar "H1"%string);(PVar "T2"%string);(PVar "H2"%string);(PVar "M"%string);(PCons (PVar "H3"%string) (PVar "T3"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("umerge3_21_3"%string, 6)) [(EVar "T1"%string);(EVar "H1"%string);(EVar "T2"%string);(EVar "H2"%string);(ECons (EVar "H3"%string) (EVar "M"%string));(EVar "T3"%string)]));([(PVar "T1"%string);(PVar "H1"%string);(PVar "T2"%string);(PVar "H2"%string);(PVar "M"%string);PNil], (ELit (Atom "true"%string)), (EApp (EFunId ("umerge2_2"%string, 4)) [(EVar "T1"%string);(EVar "T2"%string);(ECons (EVar "H2"%string) (EVar "M"%string));(EVar "H1"%string)]));([(PVar "_11"%string);(PVar "_10"%string);(PVar "_9"%string);(PVar "_8"%string);(PVar "_7"%string);(PVar "_6"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_11"%string);(EVar "_10"%string);(EVar "_9"%string);(EVar "_8"%string);(EVar "_7"%string);(EVar "_6"%string)])]))]) |};
          {| identifier := ("rumerge3_1"%string, 6) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string)]) [([(PCons (PVar "H1"%string) (PVar "T1"%string));(PVar "T2"%string);(PVar "H2"%string);(PVar "M"%string);(PVar "T3"%string);(PVar "H3"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "H1"%string);(EVar "H2"%string)]), (ECase (EValues [(EVar "T1"%string);(EVar "H1"%string);(EVar "T2"%string);(EVar "H2"%string);(EVar "M"%string);(EVar "T3"%string);(EVar "H3"%string)]) [([(PVar "_20"%string);(PVar "_21"%string);(PVar "_22"%string);(PVar "_23"%string);(PVar "_24"%string);(PVar "_25"%string);(PVar "_26"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "_23"%string);(EVar "_26"%string)]), (EApp (EFunId ("rumerge3_12_3"%string, 7)) [(EVar "_20"%string);(EVar "_22"%string);(EVar "_23"%string);(EVar "_24"%string);(EVar "_25"%string);(EVar "_26"%string);(EVar "_21"%string)]));([(PVar "_27"%string);(PVar "_28"%string);(PVar "_29"%string);(PVar "_30"%string);(PVar "_31"%string);(PVar "_32"%string);(PVar "_33"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rumerge3_2"%string, 7)) [(EVar "_27"%string);(EVar "_29"%string);(EVar "_30"%string);(EVar "_31"%string);(EVar "_32"%string);(EVar "_33"%string);(EVar "_28"%string)]))]));([(PCons (PVar "H1"%string) (PVar "T1"%string));(PVar "T2"%string);(PVar "H2"%string);(PVar "M"%string);(PVar "T3"%string);(PVar "H3"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "H1"%string);(EVar "H3"%string)]), (EApp (EFunId ("rumerge3_21_3"%string, 7)) [(EVar "T1"%string);(EVar "T2"%string);(EVar "H2"%string);(EVar "M"%string);(EVar "T3"%string);(EVar "H3"%string);(EVar "H1"%string)]));([(PCons (PVar "H1"%string) (PVar "T1"%string));(PVar "T2"%string);(PVar "H2"%string);(PVar "M"%string);(PVar "T3"%string);(PVar "H3"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rumerge3_1"%string, 6)) [(EVar "T1"%string);(EVar "T2"%string);(EVar "H2"%string);(ECons (EVar "H1"%string) (EVar "M"%string));(EVar "T3"%string);(EVar "H3"%string)]));([PNil;(PVar "T2"%string);(PVar "H2"%string);(PVar "M"%string);(PVar "T3"%string);(PVar "H3"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "H2"%string);(EVar "H3"%string)]), (EApp (EFunId ("rumerge2_2"%string, 5)) [(EVar "T2"%string);(EVar "T3"%string);(EVar "M"%string);(EVar "H3"%string);(EVar "H2"%string)]));([PNil;(PVar "T2"%string);(PVar "H2"%string);(PVar "M"%string);(PVar "T3"%string);(PVar "H3"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rumerge2_1"%string, 4)) [(EVar "T2"%string);(EVar "T3"%string);(ECons (EVar "H2"%string) (EVar "M"%string));(EVar "H3"%string)]));([(PVar "_11"%string);(PVar "_10"%string);(PVar "_9"%string);(PVar "_8"%string);(PVar "_7"%string);(PVar "_6"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_11"%string);(EVar "_10"%string);(EVar "_9"%string);(EVar "_8"%string);(EVar "_7"%string);(EVar "_6"%string)])]))]) |};
          {| identifier := ("rumerge3_12a"%string, 7) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string;"_6"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string);(EVar "_6"%string)]) [([(PVar "T1"%string);(PVar "H1"%string);(PVar "T2"%string);(PVar "H2"%string);(PVar "M"%string);(PVar "T3"%string);(PVar "H3"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "H2"%string);(EVar "H3"%string)]), (EApp (EFunId ("rumerge3_12_3"%string, 7)) [(EVar "T1"%string);(EVar "T2"%string);(EVar "H2"%string);(EVar "M"%string);(EVar "T3"%string);(EVar "H3"%string);(EVar "H1"%string)]));([(PVar "T1"%string);(PVar "H1"%string);(PVar "T2"%string);(PVar "H2"%string);(PVar "M"%string);(PVar "T3"%string);(PVar "H3"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rumerge3_2"%string, 7)) [(EVar "T1"%string);(EVar "T2"%string);(EVar "H2"%string);(EVar "M"%string);(EVar "T3"%string);(EVar "H3"%string);(EVar "H1"%string)]))]) |};
          {| identifier := ("rumerge3_2"%string, 7) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string;"_6"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string);(EVar "_6"%string)]) [([(PVar "T1"%string);(PCons (PVar "H2"%string) (PVar "T2"%string));(PVar "H2M"%string);(PVar "M"%string);(PVar "T3"%string);(PVar "H3"%string);(PVar "H1"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "H1"%string);(EVar "H2"%string)]), (ECase (EValues [(EVar "T1"%string);(EVar "H1"%string);(EVar "T2"%string);(EVar "H2"%string);(EVar "M"%string);(EVar "T3"%string);(EVar "H3"%string);(EVar "H2M"%string)]) [([(PVar "_23"%string);(PVar "_24"%string);(PVar "_25"%string);(PVar "_26"%string);(PVar "_27"%string);(PVar "_28"%string);(PVar "_29"%string);(PVar "_30"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "_26"%string);(EVar "_29"%string)]), (EApp (EFunId ("rumerge3_12_3"%string, 7)) [(EVar "_23"%string);(EVar "_25"%string);(EVar "_26"%string);(ECons (EVar "_30"%string) (EVar "_27"%string));(EVar "_28"%string);(EVar "_29"%string);(EVar "_24"%string)]));([(PVar "_31"%string);(PVar "_32"%string);(PVar "_33"%string);(PVar "_34"%string);(PVar "_35"%string);(PVar "_36"%string);(PVar "_37"%string);(PVar "_38"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rumerge3_2"%string, 7)) [(EVar "_31"%string);(EVar "_33"%string);(EVar "_34"%string);(ECons (EVar "_38"%string) (EVar "_35"%string));(EVar "_36"%string);(EVar "_37"%string);(EVar "_32"%string)]))]));([(PVar "T1"%string);(PCons (PVar "H2"%string) (PVar "T2"%string));(PVar "H2M"%string);(PVar "M"%string);(PVar "T3"%string);(PVar "H3"%string);(PVar "H1"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "H1"%string);(EVar "H2M"%string)]), (EApp (EFunId ("rumerge3_1"%string, 6)) [(EVar "T1"%string);(EVar "T2"%string);(EVar "H2"%string);(ECons (EVar "H1"%string) (EVar "M"%string));(EVar "T3"%string);(EVar "H3"%string)]));([(PVar "T1"%string);(PCons (PVar "H2"%string) (PVar "T2"%string));(PVar "H2M"%string);(PVar "M"%string);(PVar "T3"%string);(PVar "H3"%string);(PVar "H1"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "H1"%string);(EVar "H3"%string)]), (EApp (EFunId ("rumerge3_21_3"%string, 7)) [(EVar "T1"%string);(EVar "T2"%string);(EVar "H2"%string);(ECons (EVar "H2M"%string) (EVar "M"%string));(EVar "T3"%string);(EVar "H3"%string);(EVar "H1"%string)]));([(PVar "T1"%string);(PCons (PVar "H2"%string) (PVar "T2"%string));(PVar "H2M"%string);(PVar "M"%string);(PVar "T3"%string);(PVar "H3"%string);(PVar "H1"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rumerge3_1"%string, 6)) [(EVar "T1"%string);(EVar "T2"%string);(EVar "H2"%string);(ECons (EVar "H1"%string) (ECons (EVar "H2M"%string) (EVar "M"%string)));(EVar "T3"%string);(EVar "H3"%string)]));([(PVar "T1"%string);PNil;(PVar "H2M"%string);(PVar "M"%string);(PVar "T3"%string);(PVar "H3"%string);(PVar "H1"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "H1"%string);(EVar "H2M"%string)]), (EApp (EFunId ("rumerge2_1"%string, 4)) [(EVar "T1"%string);(EVar "T3"%string);(ECons (EVar "H1"%string) (EVar "M"%string));(EVar "H3"%string)]));([(PVar "T1"%string);PNil;(PVar "H2M"%string);(PVar "M"%string);(PVar "T3"%string);(PVar "H3"%string);(PVar "H1"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "H1"%string);(EVar "H3"%string)]), (EApp (EFunId ("rumerge2_2"%string, 5)) [(EVar "T1"%string);(EVar "T3"%string);(ECons (EVar "H2M"%string) (EVar "M"%string));(EVar "H3"%string);(EVar "H1"%string)]));([(PVar "T1"%string);PNil;(PVar "H2M"%string);(PVar "M"%string);(PVar "T3"%string);(PVar "H3"%string);(PVar "H1"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rumerge2_1"%string, 4)) [(EVar "T1"%string);(EVar "T3"%string);(ECons (EVar "H1"%string) (ECons (EVar "H2M"%string) (EVar "M"%string)));(EVar "H3"%string)]));([(PVar "_13"%string);(PVar "_12"%string);(PVar "_11"%string);(PVar "_10"%string);(PVar "_9"%string);(PVar "_8"%string);(PVar "_7"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_13"%string);(EVar "_12"%string);(EVar "_11"%string);(EVar "_10"%string);(EVar "_9"%string);(EVar "_8"%string);(EVar "_7"%string)])]))]) |};
          {| identifier := ("rumerge3_12b"%string, 8) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string;"_6"%string;"_7"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string);(EVar "_6"%string);(EVar "_7"%string)]) [([(PVar "T1"%string);(PVar "H1"%string);(PVar "T2"%string);(PVar "H2"%string);(PVar "M"%string);(PVar "T3"%string);(PVar "H3"%string);(PVar "H2M"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "H2"%string);(EVar "H3"%string)]), (EApp (EFunId ("rumerge3_12_3"%string, 7)) [(EVar "T1"%string);(EVar "T2"%string);(EVar "H2"%string);(ECons (EVar "H2M"%string) (EVar "M"%string));(EVar "T3"%string);(EVar "H3"%string);(EVar "H1"%string)]));([(PVar "T1"%string);(PVar "H1"%string);(PVar "T2"%string);(PVar "H2"%string);(PVar "M"%string);(PVar "T3"%string);(PVar "H3"%string);(PVar "H2M"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rumerge3_2"%string, 7)) [(EVar "T1"%string);(EVar "T2"%string);(EVar "H2"%string);(ECons (EVar "H2M"%string) (EVar "M"%string));(EVar "T3"%string);(EVar "H3"%string);(EVar "H1"%string)]))]) |};
          {| identifier := ("rumerge3_12_3"%string, 7) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string;"_6"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string);(EVar "_6"%string)]) [([(PVar "T1"%string);(PVar "T2"%string);(PVar "H2"%string);(PVar "M"%string);(PCons (PVar "H3"%string) (PVar "T3"%string));(PVar "H3M"%string);(PVar "H1"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "H2"%string);(EVar "H3"%string)]), (EApp (EFunId ("rumerge3_12_3"%string, 7)) [(EVar "T1"%string);(EVar "T2"%string);(EVar "H2"%string);(ECons (EVar "H3M"%string) (EVar "M"%string));(EVar "T3"%string);(EVar "H3"%string);(EVar "H1"%string)]));([(PVar "T1"%string);(PVar "T2"%string);(PVar "H2"%string);(PVar "M"%string);(PCons (PVar "H3"%string) (PVar "T3"%string));(PVar "H3M"%string);(PVar "H1"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "H2"%string);(EVar "H3M"%string)]), (EApp (EFunId ("rumerge3_2"%string, 7)) [(EVar "T1"%string);(EVar "T2"%string);(EVar "H2"%string);(EVar "M"%string);(EVar "T3"%string);(EVar "H3"%string);(EVar "H1"%string)]));([(PVar "T1"%string);(PVar "T2"%string);(PVar "H2"%string);(PVar "M"%string);(PCons (PVar "H3"%string) (PVar "T3"%string));(PVar "H3M"%string);(PVar "H1"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rumerge3_2"%string, 7)) [(EVar "T1"%string);(EVar "T2"%string);(EVar "H2"%string);(ECons (EVar "H3M"%string) (EVar "M"%string));(EVar "T3"%string);(EVar "H3"%string);(EVar "H1"%string)]));([(PVar "T1"%string);(PVar "T2"%string);(PVar "H2"%string);(PVar "M"%string);PNil;(PVar "H3M"%string);(PVar "H1"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "H2"%string);(EVar "H3M"%string)]), (EApp (EFunId ("rumerge2_2"%string, 5)) [(EVar "T1"%string);(EVar "T2"%string);(EVar "M"%string);(EVar "H2"%string);(EVar "H1"%string)]));([(PVar "T1"%string);(PVar "T2"%string);(PVar "H2"%string);(PVar "M"%string);PNil;(PVar "H3M"%string);(PVar "H1"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rumerge2_2"%string, 5)) [(EVar "T1"%string);(EVar "T2"%string);(ECons (EVar "H3M"%string) (EVar "M"%string));(EVar "H2"%string);(EVar "H1"%string)]));([(PVar "_13"%string);(PVar "_12"%string);(PVar "_11"%string);(PVar "_10"%string);(PVar "_9"%string);(PVar "_8"%string);(PVar "_7"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_13"%string);(EVar "_12"%string);(EVar "_11"%string);(EVar "_10"%string);(EVar "_9"%string);(EVar "_8"%string);(EVar "_7"%string)])]))]) |};
          {| identifier := ("rumerge3_21_3"%string, 7) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string;"_6"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string);(EVar "_6"%string)]) [([(PVar "T1"%string);(PVar "T2"%string);(PVar "H2"%string);(PVar "M"%string);(PCons (PVar "H3"%string) (PVar "T3"%string));(PVar "H3M"%string);(PVar "H1"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "H1"%string);(EVar "H3"%string)]), (EApp (EFunId ("rumerge3_21_3"%string, 7)) [(EVar "T1"%string);(EVar "T2"%string);(EVar "H2"%string);(ECons (EVar "H3M"%string) (EVar "M"%string));(EVar "T3"%string);(EVar "H3"%string);(EVar "H1"%string)]));([(PVar "T1"%string);(PVar "T2"%string);(PVar "H2"%string);(PVar "M"%string);(PCons (PVar "H3"%string) (PVar "T3"%string));(PVar "H3M"%string);(PVar "H1"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "H1"%string);(EVar "H3M"%string)]), (EApp (EFunId ("rumerge3_1"%string, 6)) [(EVar "T1"%string);(EVar "T2"%string);(EVar "H2"%string);(ECons (EVar "H1"%string) (EVar "M"%string));(EVar "T3"%string);(EVar "H3"%string)]));([(PVar "T1"%string);(PVar "T2"%string);(PVar "H2"%string);(PVar "M"%string);(PCons (PVar "H3"%string) (PVar "T3"%string));(PVar "H3M"%string);(PVar "H1"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rumerge3_1"%string, 6)) [(EVar "T1"%string);(EVar "T2"%string);(EVar "H2"%string);(ECons (EVar "H1"%string) (ECons (EVar "H3M"%string) (EVar "M"%string)));(EVar "T3"%string);(EVar "H3"%string)]));([(PVar "T1"%string);(PVar "T2"%string);(PVar "H2"%string);(PVar "M"%string);PNil;(PVar "H3M"%string);(PVar "H1"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "H1"%string);(EVar "H3M"%string)]), (EApp (EFunId ("rumerge2_1"%string, 4)) [(EVar "T1"%string);(EVar "T2"%string);(ECons (EVar "H1"%string) (EVar "M"%string));(EVar "H2"%string)]));([(PVar "T1"%string);(PVar "T2"%string);(PVar "H2"%string);(PVar "M"%string);PNil;(PVar "H3M"%string);(PVar "H1"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rumerge2_1"%string, 4)) [(EVar "T1"%string);(EVar "T2"%string);(ECons (EVar "H1"%string) (ECons (EVar "H3M"%string) (EVar "M"%string)));(EVar "H2"%string)]));([(PVar "_13"%string);(PVar "_12"%string);(PVar "_11"%string);(PVar "_10"%string);(PVar "_9"%string);(PVar "_8"%string);(PVar "_7"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_13"%string);(EVar "_12"%string);(EVar "_11"%string);(EVar "_10"%string);(EVar "_9"%string);(EVar "_8"%string);(EVar "_7"%string)])]))]) |};
          {| identifier := ("umerge2_1"%string, 5) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string)]) [([(PCons (PVar "H1"%string) (PVar "T1"%string));(PVar "T2"%string);(PVar "M"%string);(PVar "_HdM"%string);(PVar "H2"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "H1"%string);(EVar "H2"%string)]), (EApp (EFunId ("umerge2_1"%string, 5)) [(EVar "T1"%string);(EVar "T2"%string);(ECons (EVar "H1"%string) (EVar "M"%string));(EVar "H1"%string);(EVar "H2"%string)]));([(PCons (PVar "H1"%string) (PVar "T1"%string));(PVar "T2"%string);(PVar "M"%string);(PVar "HdM"%string);(PVar "H2"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "H2"%string);(EVar "HdM"%string)]), (EApp (EFunId ("umerge2_2"%string, 4)) [(EVar "T1"%string);(EVar "T2"%string);(EVar "M"%string);(EVar "H1"%string)]));([(PCons (PVar "H1"%string) (PVar "T1"%string));(PVar "T2"%string);(PVar "M"%string);(PVar "_HdM"%string);(PVar "H2"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("umerge2_2"%string, 4)) [(EVar "T1"%string);(EVar "T2"%string);(ECons (EVar "H2"%string) (EVar "M"%string));(EVar "H1"%string)]));([PNil;(PVar "T2"%string);(PVar "M"%string);(PVar "HdM"%string);(PVar "H2"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "H2"%string);(EVar "HdM"%string)]), (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "T2"%string);(EVar "M"%string)]));([PNil;(PVar "T2"%string);(PVar "M"%string);(PVar "_HdM"%string);(PVar "H2"%string)], (ELit (Atom "true"%string)), (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "T2"%string);(ECons (EVar "H2"%string) (EVar "M"%string))]));([(PVar "_9"%string);(PVar "_8"%string);(PVar "_7"%string);(PVar "_6"%string);(PVar "_5"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_9"%string);(EVar "_8"%string);(EVar "_7"%string);(EVar "_6"%string);(EVar "_5"%string)])]))]) |};
          {| identifier := ("umerge2_2"%string, 4) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string)]) [([(PVar "T1"%string);(PCons (PVar "H2"%string) (PVar "T2"%string));(PVar "M"%string);(PVar "H1"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "H1"%string);(EVar "H2"%string)]), (EApp (EFunId ("umerge2_1"%string, 5)) [(EVar "T1"%string);(EVar "T2"%string);(ECons (EVar "H1"%string) (EVar "M"%string));(EVar "H1"%string);(EVar "H2"%string)]));([(PVar "T1"%string);(PCons (PVar "H2"%string) (PVar "T2"%string));(PVar "M"%string);(PVar "H1"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("umerge2_2"%string, 4)) [(EVar "T1"%string);(EVar "T2"%string);(ECons (EVar "H2"%string) (EVar "M"%string));(EVar "H1"%string)]));([(PVar "T1"%string);PNil;(PVar "M"%string);(PVar "H1"%string)], (ELit (Atom "true"%string)), (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "T1"%string);(ECons (EVar "H1"%string) (EVar "M"%string))]));([(PVar "_7"%string);(PVar "_6"%string);(PVar "_5"%string);(PVar "_4"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_7"%string);(EVar "_6"%string);(EVar "_5"%string);(EVar "_4"%string)])]))]) |};
          {| identifier := ("rumerge2_1"%string, 4) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string)]) [([(PCons (PVar "H1"%string) (PVar "T1"%string));(PVar "T2"%string);(PVar "M"%string);(PVar "H2"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "H1"%string);(EVar "H2"%string)]), (EApp (EFunId ("rumerge2_2"%string, 5)) [(EVar "T1"%string);(EVar "T2"%string);(EVar "M"%string);(EVar "H2"%string);(EVar "H1"%string)]));([(PCons (PVar "H1"%string) (PVar "T1"%string));(PVar "T2"%string);(PVar "M"%string);(PVar "H2"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rumerge2_1"%string, 4)) [(EVar "T1"%string);(EVar "T2"%string);(ECons (EVar "H1"%string) (EVar "M"%string));(EVar "H2"%string)]));([PNil;(PVar "T2"%string);(PVar "M"%string);(PVar "H2"%string)], (ELit (Atom "true"%string)), (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "T2"%string);(ECons (EVar "H2"%string) (EVar "M"%string))]));([(PVar "_7"%string);(PVar "_6"%string);(PVar "_5"%string);(PVar "_4"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_7"%string);(EVar "_6"%string);(EVar "_5"%string);(EVar "_4"%string)])]))]) |};
          {| identifier := ("rumerge2_2"%string, 5) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string)]) [([(PVar "T1"%string);(PCons (PVar "H2"%string) (PVar "T2"%string));(PVar "M"%string);(PVar "H2M"%string);(PVar "H1"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "H1"%string);(EVar "H2"%string)]), (EApp (EFunId ("rumerge2_2"%string, 5)) [(EVar "T1"%string);(EVar "T2"%string);(ECons (EVar "H2M"%string) (EVar "M"%string));(EVar "H2"%string);(EVar "H1"%string)]));([(PVar "T1"%string);(PCons (PVar "H2"%string) (PVar "T2"%string));(PVar "M"%string);(PVar "H2M"%string);(PVar "H1"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "H1"%string);(EVar "H2M"%string)]), (EApp (EFunId ("rumerge2_1"%string, 4)) [(EVar "T1"%string);(EVar "T2"%string);(ECons (EVar "H1"%string) (EVar "M"%string));(EVar "H2"%string)]));([(PVar "T1"%string);(PCons (PVar "H2"%string) (PVar "T2"%string));(PVar "M"%string);(PVar "H2M"%string);(PVar "H1"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rumerge2_1"%string, 4)) [(EVar "T1"%string);(EVar "T2"%string);(ECons (EVar "H1"%string) (ECons (EVar "H2M"%string) (EVar "M"%string)));(EVar "H2"%string)]));([(PVar "T1"%string);PNil;(PVar "M"%string);(PVar "H2M"%string);(PVar "H1"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "H1"%string);(EVar "H2M"%string)]), (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "T1"%string);(ECons (EVar "H1"%string) (EVar "M"%string))]));([(PVar "T1"%string);PNil;(PVar "M"%string);(PVar "H2M"%string);(PVar "H1"%string)], (ELit (Atom "true"%string)), (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "T1"%string);(ECons (EVar "H1"%string) (ECons (EVar "H2M"%string) (EVar "M"%string)))]));([(PVar "_9"%string);(PVar "_8"%string);(PVar "_7"%string);(PVar "_6"%string);(PVar "_5"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_9"%string);(EVar "_8"%string);(EVar "_7"%string);(EVar "_6"%string);(EVar "_5"%string)])]))]) |};
          {| identifier := ("keysplit_1"%string, 8) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string;"_6"%string;"_7"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string);(EVar "_6"%string);(EVar "_7"%string)]) [([(PVar "I"%string);(PVar "X"%string);(PVar "EX"%string);(PVar "Y"%string);(PVar "EY"%string);(PCons (PVar "Z"%string) (PVar "L"%string));(PVar "R"%string);(PVar "Rs"%string)], (ELit (Atom "true"%string)), (ECase (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "I"%string);(EVar "Z"%string)]) [([(PVar "EZ"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "EY"%string);(EVar "EZ"%string)]), (EApp (EFunId ("keysplit_1"%string, 8)) [(EVar "I"%string);(EVar "Y"%string);(EVar "EY"%string);(EVar "Z"%string);(EVar "EZ"%string);(EVar "L"%string);(ECons (EVar "X"%string) (EVar "R"%string));(EVar "Rs"%string)]));([(PVar "EZ"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "EX"%string);(EVar "EZ"%string)]), (EApp (EFunId ("keysplit_1"%string, 8)) [(EVar "I"%string);(EVar "Z"%string);(EVar "EZ"%string);(EVar "Y"%string);(EVar "EY"%string);(EVar "L"%string);(ECons (EVar "X"%string) (EVar "R"%string));(EVar "Rs"%string)]));([(PVar "_EZ"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "R"%string);ENil]), (EApp (EFunId ("keysplit_1"%string, 8)) [(EVar "I"%string);(EVar "X"%string);(EVar "EX"%string);(EVar "Y"%string);(EVar "EY"%string);(EVar "L"%string);(ECons (EVar "Z"%string) ENil);(EVar "Rs"%string)]));([(PVar "EZ"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("keysplit_1_1"%string, 10)) [(EVar "I"%string);(EVar "X"%string);(EVar "EX"%string);(EVar "Y"%string);(EVar "EY"%string);(EVar "EZ"%string);(EVar "R"%string);(EVar "Rs"%string);(EVar "Z"%string);(EVar "L"%string)]))]));([(PVar "I"%string);(PVar "X"%string);(PVar "_EX"%string);(PVar "Y"%string);(PVar "_EY"%string);PNil;(PVar "R"%string);(PVar "Rs"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rkeymergel"%string, 4)) [(EVar "I"%string);(ECons (ECons (EVar "Y"%string) (ECons (EVar "X"%string) (EVar "R"%string))) (EVar "Rs"%string));ENil;(ELit (Atom "asc"%string))]));([(PVar "_16"%string);(PVar "_15"%string);(PVar "_14"%string);(PVar "_13"%string);(PVar "_12"%string);(PVar "_11"%string);(PVar "_10"%string);(PVar "_9"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_16"%string);(EVar "_15"%string);(EVar "_14"%string);(EVar "_13"%string);(EVar "_12"%string);(EVar "_11"%string);(EVar "_10"%string);(EVar "_9"%string)])]))]) |};
          {| identifier := ("keysplit_1_1"%string, 10) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string;"_6"%string;"_7"%string;"_8"%string;"_9"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string);(EVar "_6"%string);(EVar "_7"%string);(EVar "_8"%string);(EVar "_9"%string)]) [([(PVar "I"%string);(PVar "X"%string);(PVar "EX"%string);(PVar "Y"%string);(PVar "EY"%string);(PVar "ES"%string);(PVar "R"%string);(PVar "Rs"%string);(PVar "S"%string);(PCons (PVar "Z"%string) (PVar "L"%string))], (ELit (Atom "true"%string)), (ECase (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "I"%string);(EVar "Z"%string)]) [([(PVar "EZ"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "EY"%string);(EVar "EZ"%string)]), (EApp (EFunId ("keysplit_1_1"%string, 10)) [(EVar "I"%string);(EVar "Y"%string);(EVar "EY"%string);(EVar "Z"%string);(EVar "EZ"%string);(EVar "ES"%string);(ECons (EVar "X"%string) (EVar "R"%string));(EVar "Rs"%string);(EVar "S"%string);(EVar "L"%string)]));([(PVar "EZ"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "EX"%string);(EVar "EZ"%string)]), (EApp (EFunId ("keysplit_1_1"%string, 10)) [(EVar "I"%string);(EVar "Z"%string);(EVar "EZ"%string);(EVar "Y"%string);(EVar "EY"%string);(EVar "ES"%string);(ECons (EVar "X"%string) (EVar "R"%string));(EVar "Rs"%string);(EVar "S"%string);(EVar "L"%string)]));([(PVar "EZ"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "ES"%string);(EVar "EZ"%string)]), (EApp (EFunId ("keysplit_1"%string, 8)) [(EVar "I"%string);(EVar "S"%string);(EVar "ES"%string);(EVar "Z"%string);(EVar "EZ"%string);(EVar "L"%string);ENil;(ECons (ECons (EVar "Y"%string) (ECons (EVar "X"%string) (EVar "R"%string))) (EVar "Rs"%string))]));([(PVar "EZ"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("keysplit_1"%string, 8)) [(EVar "I"%string);(EVar "Z"%string);(EVar "EZ"%string);(EVar "S"%string);(EVar "ES"%string);(EVar "L"%string);ENil;(ECons (ECons (EVar "Y"%string) (ECons (EVar "X"%string) (EVar "R"%string))) (EVar "Rs"%string))]))]));([(PVar "I"%string);(PVar "X"%string);(PVar "_EX"%string);(PVar "Y"%string);(PVar "_EY"%string);(PVar "_ES"%string);(PVar "R"%string);(PVar "Rs"%string);(PVar "S"%string);PNil], (ELit (Atom "true"%string)), (EApp (EFunId ("rkeymergel"%string, 4)) [(EVar "I"%string);(ECons (ECons (EVar "S"%string) ENil) (ECons (ECons (EVar "Y"%string) (ECons (EVar "X"%string) (EVar "R"%string))) (EVar "Rs"%string)));ENil;(ELit (Atom "asc"%string))]));([(PVar "_20"%string);(PVar "_19"%string);(PVar "_18"%string);(PVar "_17"%string);(PVar "_16"%string);(PVar "_15"%string);(PVar "_14"%string);(PVar "_13"%string);(PVar "_12"%string);(PVar "_11"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_20"%string);(EVar "_19"%string);(EVar "_18"%string);(EVar "_17"%string);(EVar "_16"%string);(EVar "_15"%string);(EVar "_14"%string);(EVar "_13"%string);(EVar "_12"%string);(EVar "_11"%string)])]))]) |};
          {| identifier := ("keysplit_2"%string, 8) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string;"_6"%string;"_7"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string);(EVar "_6"%string);(EVar "_7"%string)]) [([(PVar "I"%string);(PVar "X"%string);(PVar "EX"%string);(PVar "Y"%string);(PVar "EY"%string);(PCons (PVar "Z"%string) (PVar "L"%string));(PVar "R"%string);(PVar "Rs"%string)], (ELit (Atom "true"%string)), (ECase (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "I"%string);(EVar "Z"%string)]) [([(PVar "EZ"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom ">"%string)) [(EVar "EY"%string);(EVar "EZ"%string)]), (EApp (EFunId ("keysplit_2"%string, 8)) [(EVar "I"%string);(EVar "Y"%string);(EVar "EY"%string);(EVar "Z"%string);(EVar "EZ"%string);(EVar "L"%string);(ECons (EVar "X"%string) (EVar "R"%string));(EVar "Rs"%string)]));([(PVar "EZ"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom ">"%string)) [(EVar "EX"%string);(EVar "EZ"%string)]), (EApp (EFunId ("keysplit_2"%string, 8)) [(EVar "I"%string);(EVar "Z"%string);(EVar "EZ"%string);(EVar "Y"%string);(EVar "EY"%string);(EVar "L"%string);(ECons (EVar "X"%string) (EVar "R"%string));(EVar "Rs"%string)]));([(PVar "_EZ"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "R"%string);ENil]), (EApp (EFunId ("keysplit_2"%string, 8)) [(EVar "I"%string);(EVar "X"%string);(EVar "EX"%string);(EVar "Y"%string);(EVar "EY"%string);(EVar "L"%string);(ECons (EVar "Z"%string) ENil);(EVar "Rs"%string)]));([(PVar "EZ"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("keysplit_2_1"%string, 10)) [(EVar "I"%string);(EVar "X"%string);(EVar "EX"%string);(EVar "Y"%string);(EVar "EY"%string);(EVar "EZ"%string);(EVar "R"%string);(EVar "Rs"%string);(EVar "Z"%string);(EVar "L"%string)]))]));([(PVar "I"%string);(PVar "X"%string);(PVar "_EX"%string);(PVar "Y"%string);(PVar "_EY"%string);PNil;(PVar "R"%string);(PVar "Rs"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("keymergel"%string, 4)) [(EVar "I"%string);(ECons (ECons (EVar "Y"%string) (ECons (EVar "X"%string) (EVar "R"%string))) (EVar "Rs"%string));ENil;(ELit (Atom "desc"%string))]));([(PVar "_16"%string);(PVar "_15"%string);(PVar "_14"%string);(PVar "_13"%string);(PVar "_12"%string);(PVar "_11"%string);(PVar "_10"%string);(PVar "_9"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_16"%string);(EVar "_15"%string);(EVar "_14"%string);(EVar "_13"%string);(EVar "_12"%string);(EVar "_11"%string);(EVar "_10"%string);(EVar "_9"%string)])]))]) |};
          {| identifier := ("keysplit_2_1"%string, 10) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string;"_6"%string;"_7"%string;"_8"%string;"_9"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string);(EVar "_6"%string);(EVar "_7"%string);(EVar "_8"%string);(EVar "_9"%string)]) [([(PVar "I"%string);(PVar "X"%string);(PVar "EX"%string);(PVar "Y"%string);(PVar "EY"%string);(PVar "ES"%string);(PVar "R"%string);(PVar "Rs"%string);(PVar "S"%string);(PCons (PVar "Z"%string) (PVar "L"%string))], (ELit (Atom "true"%string)), (ECase (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "I"%string);(EVar "Z"%string)]) [([(PVar "EZ"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom ">"%string)) [(EVar "EY"%string);(EVar "EZ"%string)]), (EApp (EFunId ("keysplit_2_1"%string, 10)) [(EVar "I"%string);(EVar "Y"%string);(EVar "EY"%string);(EVar "Z"%string);(EVar "EZ"%string);(EVar "ES"%string);(ECons (EVar "X"%string) (EVar "R"%string));(EVar "Rs"%string);(EVar "S"%string);(EVar "L"%string)]));([(PVar "EZ"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom ">"%string)) [(EVar "EX"%string);(EVar "EZ"%string)]), (EApp (EFunId ("keysplit_2_1"%string, 10)) [(EVar "I"%string);(EVar "Z"%string);(EVar "EZ"%string);(EVar "Y"%string);(EVar "EY"%string);(EVar "ES"%string);(ECons (EVar "X"%string) (EVar "R"%string));(EVar "Rs"%string);(EVar "S"%string);(EVar "L"%string)]));([(PVar "EZ"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom ">"%string)) [(EVar "ES"%string);(EVar "EZ"%string)]), (EApp (EFunId ("keysplit_2"%string, 8)) [(EVar "I"%string);(EVar "S"%string);(EVar "ES"%string);(EVar "Z"%string);(EVar "EZ"%string);(EVar "L"%string);ENil;(ECons (ECons (EVar "Y"%string) (ECons (EVar "X"%string) (EVar "R"%string))) (EVar "Rs"%string))]));([(PVar "EZ"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("keysplit_2"%string, 8)) [(EVar "I"%string);(EVar "Z"%string);(EVar "EZ"%string);(EVar "S"%string);(EVar "ES"%string);(EVar "L"%string);ENil;(ECons (ECons (EVar "Y"%string) (ECons (EVar "X"%string) (EVar "R"%string))) (EVar "Rs"%string))]))]));([(PVar "I"%string);(PVar "X"%string);(PVar "_EX"%string);(PVar "Y"%string);(PVar "_EY"%string);(PVar "_ES"%string);(PVar "R"%string);(PVar "Rs"%string);(PVar "S"%string);PNil], (ELit (Atom "true"%string)), (EApp (EFunId ("keymergel"%string, 4)) [(EVar "I"%string);(ECons (ECons (EVar "S"%string) ENil) (ECons (ECons (EVar "Y"%string) (ECons (EVar "X"%string) (EVar "R"%string))) (EVar "Rs"%string)));ENil;(ELit (Atom "desc"%string))]));([(PVar "_20"%string);(PVar "_19"%string);(PVar "_18"%string);(PVar "_17"%string);(PVar "_16"%string);(PVar "_15"%string);(PVar "_14"%string);(PVar "_13"%string);(PVar "_12"%string);(PVar "_11"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_20"%string);(EVar "_19"%string);(EVar "_18"%string);(EVar "_17"%string);(EVar "_16"%string);(EVar "_15"%string);(EVar "_14"%string);(EVar "_13"%string);(EVar "_12"%string);(EVar "_11"%string)])]))]) |};
          {| identifier := ("keymergel"%string, 4) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string)]) [([(PVar "I"%string);(PCons (PVar "T1"%string) (PCons (PCons (PVar "H2"%string) (PVar "T2"%string)) (PCons (PCons (PVar "H3"%string) (PVar "T3"%string)) (PVar "L"%string))));(PVar "Acc"%string);(PVar "O"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "O"%string);(ELit (Atom "asc"%string))]), (ELet ["_5"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "I"%string);(EVar "H2"%string)]) (ELet ["_4"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "I"%string);(EVar "H3"%string)]) (ELet ["M"%string] (EApp (EFunId ("keymerge3_1"%string, 10)) [(EVar "I"%string);(EVar "T1"%string);ENil;(EVar "O"%string);(EVar "_5"%string);(EVar "H2"%string);(EVar "T2"%string);(EVar "_4"%string);(EVar "H3"%string);(EVar "T3"%string)]) (EApp (EFunId ("keymergel"%string, 4)) [(EVar "I"%string);(EVar "L"%string);(ECons (EVar "M"%string) (EVar "Acc"%string));(EVar "O"%string)])))));([(PVar "I"%string);(PCons (PCons (PVar "H3"%string) (PVar "T3"%string)) (PCons (PCons (PVar "H2"%string) (PVar "T2"%string)) (PCons (PVar "T1"%string) (PVar "L"%string))));(PVar "Acc"%string);(PVar "O"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "O"%string);(ELit (Atom "desc"%string))]), (ELet ["_8"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "I"%string);(EVar "H2"%string)]) (ELet ["_7"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "I"%string);(EVar "H3"%string)]) (ELet ["M"%string] (EApp (EFunId ("keymerge3_1"%string, 10)) [(EVar "I"%string);(EVar "T1"%string);ENil;(EVar "O"%string);(EVar "_8"%string);(EVar "H2"%string);(EVar "T2"%string);(EVar "_7"%string);(EVar "H3"%string);(EVar "T3"%string)]) (EApp (EFunId ("keymergel"%string, 4)) [(EVar "I"%string);(EVar "L"%string);(ECons (EVar "M"%string) (EVar "Acc"%string));(EVar "O"%string)])))));([(PVar "I"%string);(PCons (PVar "T1"%string) (PCons (PCons (PVar "H2"%string) (PVar "T2"%string)) (PVar "L"%string)));(PVar "Acc"%string);(PLit (Atom "asc"%string))], (ELit (Atom "true"%string)), (ELet ["_10"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "I"%string);(EVar "H2"%string)]) (ELet ["_11"%string] (EApp (EFunId ("keymerge2_1"%string, 6)) [(EVar "I"%string);(EVar "T1"%string);(EVar "_10"%string);(EVar "H2"%string);(EVar "T2"%string);ENil]) (EApp (EFunId ("keymergel"%string, 4)) [(EVar "I"%string);(EVar "L"%string);(ECons (EVar "_11"%string) (EVar "Acc"%string));(ELit (Atom "asc"%string))]))));([(PVar "I"%string);(PCons (PCons (PVar "H2"%string) (PVar "T2"%string)) (PCons (PVar "T1"%string) (PVar "L"%string)));(PVar "Acc"%string);(PLit (Atom "desc"%string))], (ELit (Atom "true"%string)), (ELet ["_12"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "I"%string);(EVar "H2"%string)]) (ELet ["_13"%string] (EApp (EFunId ("keymerge2_1"%string, 6)) [(EVar "I"%string);(EVar "T1"%string);(EVar "_12"%string);(EVar "H2"%string);(EVar "T2"%string);ENil]) (EApp (EFunId ("keymergel"%string, 4)) [(EVar "I"%string);(EVar "L"%string);(ECons (EVar "_13"%string) (EVar "Acc"%string));(ELit (Atom "desc"%string))]))));([(PVar "_I"%string);(PCons (PVar "L"%string) PNil);PNil;(PVar "_O"%string)], (ELit (Atom "true"%string)), (EVar "L"%string));([(PVar "I"%string);(PCons (PVar "L"%string) PNil);(PVar "Acc"%string);(PVar "O"%string)], (ELit (Atom "true"%string)), (ELet ["_14"%string] (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "L"%string);ENil]) (EApp (EFunId ("rkeymergel"%string, 4)) [(EVar "I"%string);(ECons (EVar "_14"%string) (EVar "Acc"%string));ENil;(EVar "O"%string)])));([(PVar "I"%string);PNil;(PVar "Acc"%string);(PVar "O"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rkeymergel"%string, 4)) [(EVar "I"%string);(EVar "Acc"%string);ENil;(EVar "O"%string)]));([(PVar "_18"%string);(PVar "_17"%string);(PVar "_16"%string);(PVar "_15"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_18"%string);(EVar "_17"%string);(EVar "_16"%string);(EVar "_15"%string)])]))]) |};
          {| identifier := ("rkeymergel"%string, 4) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string)]) [([(PVar "I"%string);(PCons (PCons (PVar "H3"%string) (PVar "T3"%string)) (PCons (PCons (PVar "H2"%string) (PVar "T2"%string)) (PCons (PVar "T1"%string) (PVar "L"%string))));(PVar "Acc"%string);(PVar "O"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "O"%string);(ELit (Atom "asc"%string))]), (ELet ["_5"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "I"%string);(EVar "H2"%string)]) (ELet ["_4"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "I"%string);(EVar "H3"%string)]) (ELet ["M"%string] (EApp (EFunId ("rkeymerge3_1"%string, 10)) [(EVar "I"%string);(EVar "T1"%string);ENil;(EVar "O"%string);(EVar "_5"%string);(EVar "H2"%string);(EVar "T2"%string);(EVar "_4"%string);(EVar "H3"%string);(EVar "T3"%string)]) (EApp (EFunId ("rkeymergel"%string, 4)) [(EVar "I"%string);(EVar "L"%string);(ECons (EVar "M"%string) (EVar "Acc"%string));(EVar "O"%string)])))));([(PVar "I"%string);(PCons (PVar "T1"%string) (PCons (PCons (PVar "H2"%string) (PVar "T2"%string)) (PCons (PCons (PVar "H3"%string) (PVar "T3"%string)) (PVar "L"%string))));(PVar "Acc"%string);(PVar "O"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "O"%string);(ELit (Atom "desc"%string))]), (ELet ["_8"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "I"%string);(EVar "H2"%string)]) (ELet ["_7"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "I"%string);(EVar "H3"%string)]) (ELet ["M"%string] (EApp (EFunId ("rkeymerge3_1"%string, 10)) [(EVar "I"%string);(EVar "T1"%string);ENil;(EVar "O"%string);(EVar "_8"%string);(EVar "H2"%string);(EVar "T2"%string);(EVar "_7"%string);(EVar "H3"%string);(EVar "T3"%string)]) (EApp (EFunId ("rkeymergel"%string, 4)) [(EVar "I"%string);(EVar "L"%string);(ECons (EVar "M"%string) (EVar "Acc"%string));(EVar "O"%string)])))));([(PVar "I"%string);(PCons (PCons (PVar "H2"%string) (PVar "T2"%string)) (PCons (PVar "T1"%string) (PVar "L"%string)));(PVar "Acc"%string);(PLit (Atom "asc"%string))], (ELit (Atom "true"%string)), (ELet ["_10"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "I"%string);(EVar "H2"%string)]) (ELet ["_11"%string] (EApp (EFunId ("rkeymerge2_1"%string, 6)) [(EVar "I"%string);(EVar "T1"%string);(EVar "_10"%string);(EVar "H2"%string);(EVar "T2"%string);ENil]) (EApp (EFunId ("rkeymergel"%string, 4)) [(EVar "I"%string);(EVar "L"%string);(ECons (EVar "_11"%string) (EVar "Acc"%string));(ELit (Atom "asc"%string))]))));([(PVar "I"%string);(PCons (PVar "T1"%string) (PCons (PCons (PVar "H2"%string) (PVar "T2"%string)) (PVar "L"%string)));(PVar "Acc"%string);(PLit (Atom "desc"%string))], (ELit (Atom "true"%string)), (ELet ["_12"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "I"%string);(EVar "H2"%string)]) (ELet ["_13"%string] (EApp (EFunId ("rkeymerge2_1"%string, 6)) [(EVar "I"%string);(EVar "T1"%string);(EVar "_12"%string);(EVar "H2"%string);(EVar "T2"%string);ENil]) (EApp (EFunId ("rkeymergel"%string, 4)) [(EVar "I"%string);(EVar "L"%string);(ECons (EVar "_13"%string) (EVar "Acc"%string));(ELit (Atom "desc"%string))]))));([(PVar "I"%string);(PCons (PVar "L"%string) PNil);(PVar "Acc"%string);(PVar "O"%string)], (ELit (Atom "true"%string)), (ELet ["_14"%string] (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "L"%string);ENil]) (EApp (EFunId ("keymergel"%string, 4)) [(EVar "I"%string);(ECons (EVar "_14"%string) (EVar "Acc"%string));ENil;(EVar "O"%string)])));([(PVar "I"%string);PNil;(PVar "Acc"%string);(PVar "O"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("keymergel"%string, 4)) [(EVar "I"%string);(EVar "Acc"%string);ENil;(EVar "O"%string)]));([(PVar "_18"%string);(PVar "_17"%string);(PVar "_16"%string);(PVar "_15"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_18"%string);(EVar "_17"%string);(EVar "_16"%string);(EVar "_15"%string)])]))]) |};
          {| identifier := ("keymerge3_1"%string, 10) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string;"_6"%string;"_7"%string;"_8"%string;"_9"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string);(EVar "_6"%string);(EVar "_7"%string);(EVar "_8"%string);(EVar "_9"%string)]) [([(PVar "I"%string);(PCons (PVar "H1"%string) (PVar "T1"%string));(PVar "M"%string);(PVar "D"%string);(PVar "E2"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "E3"%string);(PVar "H3"%string);(PVar "T3"%string)], (ELit (Atom "true"%string)), (ECase (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "I"%string);(EVar "H1"%string)]) [([(PVar "E1"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "E1"%string);(EVar "E2"%string)]), (ECase (EValues [(EVar "I"%string);(EVar "E1"%string);(EVar "H1"%string);(EVar "T1"%string);(EVar "E2"%string);(EVar "H2"%string);(EVar "T2"%string);(EVar "E3"%string);(EVar "H3"%string);(EVar "T3"%string);(EVar "M"%string);(EVar "D"%string)]) [([(PVar "_34"%string);(PVar "_35"%string);(PVar "_36"%string);(PVar "_37"%string);(PVar "_38"%string);(PVar "_39"%string);(PVar "_40"%string);(PVar "_41"%string);(PVar "_42"%string);(PVar "_43"%string);(PVar "_44"%string);(PVar "_45"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "_35"%string);(EVar "_41"%string)]), (EApp (EFunId ("keymerge3_1"%string, 10)) [(EVar "_34"%string);(EVar "_37"%string);(ECons (EVar "_36"%string) (EVar "_44"%string));(EVar "_45"%string);(EVar "_38"%string);(EVar "_39"%string);(EVar "_40"%string);(EVar "_41"%string);(EVar "_42"%string);(EVar "_43"%string)]));([(PVar "_46"%string);(PVar "_47"%string);(PVar "_48"%string);(PVar "_49"%string);(PVar "_50"%string);(PVar "_51"%string);(PVar "_52"%string);(PVar "_E3"%string);(PVar "_53"%string);(PVar "_54"%string);(PVar "_55"%string);(PVar "_D"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("keymerge3_12_3"%string, 9)) [(EVar "_46"%string);(EVar "_47"%string);(EVar "_48"%string);(EVar "_49"%string);(EVar "_50"%string);(EVar "_51"%string);(EVar "_52"%string);(EVar "_54"%string);(ECons (EVar "_53"%string) (EVar "_55"%string))]))]));([(PVar "E1"%string)], (ELit (Atom "true"%string)), (ECase (EValues [(EVar "I"%string);(EVar "E1"%string);(EVar "H1"%string);(EVar "T1"%string);(EVar "E2"%string);(EVar "H2"%string);(EVar "T2"%string);(EVar "E3"%string);(EVar "H3"%string);(EVar "T3"%string);(EVar "M"%string);(EVar "T2"%string)]) [([(PVar "_66"%string);(PVar "_67"%string);(PVar "_68"%string);(PVar "_69"%string);(PVar "_70"%string);(PVar "_71"%string);(PVar "_72"%string);(PVar "_73"%string);(PVar "_74"%string);(PVar "_75"%string);(PVar "_76"%string);(PVar "_77"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "_70"%string);(EVar "_73"%string)]), (EApp (EFunId ("keymerge3_2"%string, 10)) [(EVar "_66"%string);(EVar "_67"%string);(EVar "_68"%string);(EVar "_69"%string);(EVar "_72"%string);(ECons (EVar "_71"%string) (EVar "_76"%string));(EVar "_77"%string);(EVar "_73"%string);(EVar "_74"%string);(EVar "_75"%string)]));([(PVar "_78"%string);(PVar "_79"%string);(PVar "_80"%string);(PVar "_81"%string);(PVar "_82"%string);(PVar "_83"%string);(PVar "_84"%string);(PVar "_E3"%string);(PVar "_85"%string);(PVar "_86"%string);(PVar "_87"%string);(PVar "_D"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("keymerge3_21_3"%string, 9)) [(EVar "_78"%string);(EVar "_79"%string);(EVar "_80"%string);(EVar "_81"%string);(EVar "_82"%string);(EVar "_83"%string);(EVar "_84"%string);(EVar "_86"%string);(ECons (EVar "_85"%string) (EVar "_87"%string))]))]))]));([(PVar "I"%string);PNil;(PVar "M"%string);(PVar "_D"%string);(PVar "E2"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "E3"%string);(PVar "H3"%string);(PVar "T3"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "E2"%string);(EVar "E3"%string)]), (EApp (EFunId ("keymerge2_1"%string, 6)) [(EVar "I"%string);(EVar "T2"%string);(EVar "E3"%string);(EVar "H3"%string);(EVar "T3"%string);(ECons (EVar "H2"%string) (EVar "M"%string))]));([(PVar "I"%string);PNil;(PVar "M"%string);(PVar "_D"%string);(PVar "E2"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "_E3"%string);(PVar "H3"%string);(PVar "T3"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("keymerge2_2"%string, 7)) [(EVar "I"%string);(EVar "T2"%string);(EVar "E2"%string);(EVar "H3"%string);(EVar "T3"%string);(EVar "M"%string);(EVar "H2"%string)]));([(PVar "_20"%string);(PVar "_19"%string);(PVar "_18"%string);(PVar "_17"%string);(PVar "_16"%string);(PVar "_15"%string);(PVar "_14"%string);(PVar "_13"%string);(PVar "_12"%string);(PVar "_11"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_20"%string);(EVar "_19"%string);(EVar "_18"%string);(EVar "_17"%string);(EVar "_16"%string);(EVar "_15"%string);(EVar "_14"%string);(EVar "_13"%string);(EVar "_12"%string);(EVar "_11"%string)])]))]) |};
          {| identifier := ("keymerge3_2"%string, 10) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string;"_6"%string;"_7"%string;"_8"%string;"_9"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string);(EVar "_6"%string);(EVar "_7"%string);(EVar "_8"%string);(EVar "_9"%string)]) [([(PVar "I"%string);(PVar "E1"%string);(PVar "H1"%string);(PVar "T1"%string);(PCons (PVar "H2"%string) (PVar "T2"%string));(PVar "M"%string);(PVar "D"%string);(PVar "E3"%string);(PVar "H3"%string);(PVar "T3"%string)], (ELit (Atom "true"%string)), (ECase (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "I"%string);(EVar "H2"%string)]) [([(PVar "E2"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "E1"%string);(EVar "E2"%string)]), (ECase (EValues [(EVar "I"%string);(EVar "E1"%string);(EVar "H1"%string);(EVar "T1"%string);(EVar "E2"%string);(EVar "H2"%string);(EVar "T2"%string);(EVar "E3"%string);(EVar "H3"%string);(EVar "T3"%string);(EVar "M"%string);(EVar "T1"%string)]) [([(PVar "_34"%string);(PVar "_35"%string);(PVar "_36"%string);(PVar "_37"%string);(PVar "_38"%string);(PVar "_39"%string);(PVar "_40"%string);(PVar "_41"%string);(PVar "_42"%string);(PVar "_43"%string);(PVar "_44"%string);(PVar "_45"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "_35"%string);(EVar "_41"%string)]), (EApp (EFunId ("keymerge3_1"%string, 10)) [(EVar "_34"%string);(EVar "_37"%string);(ECons (EVar "_36"%string) (EVar "_44"%string));(EVar "_45"%string);(EVar "_38"%string);(EVar "_39"%string);(EVar "_40"%string);(EVar "_41"%string);(EVar "_42"%string);(EVar "_43"%string)]));([(PVar "_46"%string);(PVar "_47"%string);(PVar "_48"%string);(PVar "_49"%string);(PVar "_50"%string);(PVar "_51"%string);(PVar "_52"%string);(PVar "_E3"%string);(PVar "_53"%string);(PVar "_54"%string);(PVar "_55"%string);(PVar "_D"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("keymerge3_12_3"%string, 9)) [(EVar "_46"%string);(EVar "_47"%string);(EVar "_48"%string);(EVar "_49"%string);(EVar "_50"%string);(EVar "_51"%string);(EVar "_52"%string);(EVar "_54"%string);(ECons (EVar "_53"%string) (EVar "_55"%string))]))]));([(PVar "E2"%string)], (ELit (Atom "true"%string)), (ECase (EValues [(EVar "I"%string);(EVar "E1"%string);(EVar "H1"%string);(EVar "T1"%string);(EVar "E2"%string);(EVar "H2"%string);(EVar "T2"%string);(EVar "E3"%string);(EVar "H3"%string);(EVar "T3"%string);(EVar "M"%string);(EVar "D"%string)]) [([(PVar "_66"%string);(PVar "_67"%string);(PVar "_68"%string);(PVar "_69"%string);(PVar "_70"%string);(PVar "_71"%string);(PVar "_72"%string);(PVar "_73"%string);(PVar "_74"%string);(PVar "_75"%string);(PVar "_76"%string);(PVar "_77"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "_70"%string);(EVar "_73"%string)]), (EApp (EFunId ("keymerge3_2"%string, 10)) [(EVar "_66"%string);(EVar "_67"%string);(EVar "_68"%string);(EVar "_69"%string);(EVar "_72"%string);(ECons (EVar "_71"%string) (EVar "_76"%string));(EVar "_77"%string);(EVar "_73"%string);(EVar "_74"%string);(EVar "_75"%string)]));([(PVar "_78"%string);(PVar "_79"%string);(PVar "_80"%string);(PVar "_81"%string);(PVar "_82"%string);(PVar "_83"%string);(PVar "_84"%string);(PVar "_E3"%string);(PVar "_85"%string);(PVar "_86"%string);(PVar "_87"%string);(PVar "_D"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("keymerge3_21_3"%string, 9)) [(EVar "_78"%string);(EVar "_79"%string);(EVar "_80"%string);(EVar "_81"%string);(EVar "_82"%string);(EVar "_83"%string);(EVar "_84"%string);(EVar "_86"%string);(ECons (EVar "_85"%string) (EVar "_87"%string))]))]))]));([(PVar "I"%string);(PVar "E1"%string);(PVar "H1"%string);(PVar "T1"%string);PNil;(PVar "M"%string);(PVar "_D"%string);(PVar "E3"%string);(PVar "H3"%string);(PVar "T3"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "E1"%string);(EVar "E3"%string)]), (EApp (EFunId ("keymerge2_1"%string, 6)) [(EVar "I"%string);(EVar "T1"%string);(EVar "E3"%string);(EVar "H3"%string);(EVar "T3"%string);(ECons (EVar "H1"%string) (EVar "M"%string))]));([(PVar "I"%string);(PVar "E1"%string);(PVar "H1"%string);(PVar "T1"%string);PNil;(PVar "M"%string);(PVar "_D"%string);(PVar "_E3"%string);(PVar "H3"%string);(PVar "T3"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("keymerge2_2"%string, 7)) [(EVar "I"%string);(EVar "T1"%string);(EVar "E1"%string);(EVar "H3"%string);(EVar "T3"%string);(EVar "M"%string);(EVar "H1"%string)]));([(PVar "_20"%string);(PVar "_19"%string);(PVar "_18"%string);(PVar "_17"%string);(PVar "_16"%string);(PVar "_15"%string);(PVar "_14"%string);(PVar "_13"%string);(PVar "_12"%string);(PVar "_11"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_20"%string);(EVar "_19"%string);(EVar "_18"%string);(EVar "_17"%string);(EVar "_16"%string);(EVar "_15"%string);(EVar "_14"%string);(EVar "_13"%string);(EVar "_12"%string);(EVar "_11"%string)])]))]) |};
          {| identifier := ("keymerge3_12"%string, 12) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string;"_6"%string;"_7"%string;"_8"%string;"_9"%string;"_10"%string;"_11"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string);(EVar "_6"%string);(EVar "_7"%string);(EVar "_8"%string);(EVar "_9"%string);(EVar "_10"%string);(EVar "_11"%string)]) [([(PVar "I"%string);(PVar "E1"%string);(PVar "H1"%string);(PVar "T1"%string);(PVar "E2"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "E3"%string);(PVar "H3"%string);(PVar "T3"%string);(PVar "M"%string);(PVar "D"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "E1"%string);(EVar "E3"%string)]), (EApp (EFunId ("keymerge3_1"%string, 10)) [(EVar "I"%string);(EVar "T1"%string);(ECons (EVar "H1"%string) (EVar "M"%string));(EVar "D"%string);(EVar "E2"%string);(EVar "H2"%string);(EVar "T2"%string);(EVar "E3"%string);(EVar "H3"%string);(EVar "T3"%string)]));([(PVar "I"%string);(PVar "E1"%string);(PVar "H1"%string);(PVar "T1"%string);(PVar "E2"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "_E3"%string);(PVar "H3"%string);(PVar "T3"%string);(PVar "M"%string);(PVar "_D"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("keymerge3_12_3"%string, 9)) [(EVar "I"%string);(EVar "E1"%string);(EVar "H1"%string);(EVar "T1"%string);(EVar "E2"%string);(EVar "H2"%string);(EVar "T2"%string);(EVar "T3"%string);(ECons (EVar "H3"%string) (EVar "M"%string))]))]) |};
          {| identifier := ("keymerge3_12_3"%string, 9) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string;"_6"%string;"_7"%string;"_8"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string);(EVar "_6"%string);(EVar "_7"%string);(EVar "_8"%string)]) [([(PVar "I"%string);(PVar "E1"%string);(PVar "H1"%string);(PVar "T1"%string);(PVar "E2"%string);(PVar "H2"%string);(PVar "T2"%string);(PCons (PVar "H3"%string) (PVar "T3"%string));(PVar "M"%string)], (ELit (Atom "true"%string)), (ECase (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "I"%string);(EVar "H3"%string)]) [([(PVar "E3"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "E1"%string);(EVar "E3"%string)]), (EApp (EFunId ("keymerge3_1"%string, 10)) [(EVar "I"%string);(EVar "T1"%string);(ECons (EVar "H1"%string) (EVar "M"%string));(EVar "T1"%string);(EVar "E2"%string);(EVar "H2"%string);(EVar "T2"%string);(EVar "E3"%string);(EVar "H3"%string);(EVar "T3"%string)]));([(PVar "_E3"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("keymerge3_12_3"%string, 9)) [(EVar "I"%string);(EVar "E1"%string);(EVar "H1"%string);(EVar "T1"%string);(EVar "E2"%string);(EVar "H2"%string);(EVar "T2"%string);(EVar "T3"%string);(ECons (EVar "H3"%string) (EVar "M"%string))]))]));([(PVar "I"%string);(PVar "_E1"%string);(PVar "H1"%string);(PVar "T1"%string);(PVar "E2"%string);(PVar "H2"%string);(PVar "T2"%string);PNil;(PVar "M"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("keymerge2_1"%string, 6)) [(EVar "I"%string);(EVar "T1"%string);(EVar "E2"%string);(EVar "H2"%string);(EVar "T2"%string);(ECons (EVar "H1"%string) (EVar "M"%string))]));([(PVar "_18"%string);(PVar "_17"%string);(PVar "_16"%string);(PVar "_15"%string);(PVar "_14"%string);(PVar "_13"%string);(PVar "_12"%string);(PVar "_11"%string);(PVar "_10"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_18"%string);(EVar "_17"%string);(EVar "_16"%string);(EVar "_15"%string);(EVar "_14"%string);(EVar "_13"%string);(EVar "_12"%string);(EVar "_11"%string);(EVar "_10"%string)])]))]) |};
          {| identifier := ("keymerge3_21"%string, 12) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string;"_6"%string;"_7"%string;"_8"%string;"_9"%string;"_10"%string;"_11"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string);(EVar "_6"%string);(EVar "_7"%string);(EVar "_8"%string);(EVar "_9"%string);(EVar "_10"%string);(EVar "_11"%string)]) [([(PVar "I"%string);(PVar "E1"%string);(PVar "H1"%string);(PVar "T1"%string);(PVar "E2"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "E3"%string);(PVar "H3"%string);(PVar "T3"%string);(PVar "M"%string);(PVar "D"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "E2"%string);(EVar "E3"%string)]), (EApp (EFunId ("keymerge3_2"%string, 10)) [(EVar "I"%string);(EVar "E1"%string);(EVar "H1"%string);(EVar "T1"%string);(EVar "T2"%string);(ECons (EVar "H2"%string) (EVar "M"%string));(EVar "D"%string);(EVar "E3"%string);(EVar "H3"%string);(EVar "T3"%string)]));([(PVar "I"%string);(PVar "E1"%string);(PVar "H1"%string);(PVar "T1"%string);(PVar "E2"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "_E3"%string);(PVar "H3"%string);(PVar "T3"%string);(PVar "M"%string);(PVar "_D"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("keymerge3_21_3"%string, 9)) [(EVar "I"%string);(EVar "E1"%string);(EVar "H1"%string);(EVar "T1"%string);(EVar "E2"%string);(EVar "H2"%string);(EVar "T2"%string);(EVar "T3"%string);(ECons (EVar "H3"%string) (EVar "M"%string))]))]) |};
          {| identifier := ("keymerge3_21_3"%string, 9) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string;"_6"%string;"_7"%string;"_8"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string);(EVar "_6"%string);(EVar "_7"%string);(EVar "_8"%string)]) [([(PVar "I"%string);(PVar "E1"%string);(PVar "H1"%string);(PVar "T1"%string);(PVar "E2"%string);(PVar "H2"%string);(PVar "T2"%string);(PCons (PVar "H3"%string) (PVar "T3"%string));(PVar "M"%string)], (ELit (Atom "true"%string)), (ECase (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "I"%string);(EVar "H3"%string)]) [([(PVar "E3"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "E2"%string);(EVar "E3"%string)]), (EApp (EFunId ("keymerge3_2"%string, 10)) [(EVar "I"%string);(EVar "E1"%string);(EVar "H1"%string);(EVar "T1"%string);(EVar "T2"%string);(ECons (EVar "H2"%string) (EVar "M"%string));(EVar "T2"%string);(EVar "E3"%string);(EVar "H3"%string);(EVar "T3"%string)]));([(PVar "_E3"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("keymerge3_21_3"%string, 9)) [(EVar "I"%string);(EVar "E1"%string);(EVar "H1"%string);(EVar "T1"%string);(EVar "E2"%string);(EVar "H2"%string);(EVar "T2"%string);(EVar "T3"%string);(ECons (EVar "H3"%string) (EVar "M"%string))]))]));([(PVar "I"%string);(PVar "E1"%string);(PVar "H1"%string);(PVar "T1"%string);(PVar "_E2"%string);(PVar "H2"%string);(PVar "T2"%string);PNil;(PVar "M"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("keymerge2_2"%string, 7)) [(EVar "I"%string);(EVar "T1"%string);(EVar "E1"%string);(EVar "H2"%string);(EVar "T2"%string);(EVar "M"%string);(EVar "H1"%string)]));([(PVar "_18"%string);(PVar "_17"%string);(PVar "_16"%string);(PVar "_15"%string);(PVar "_14"%string);(PVar "_13"%string);(PVar "_12"%string);(PVar "_11"%string);(PVar "_10"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_18"%string);(EVar "_17"%string);(EVar "_16"%string);(EVar "_15"%string);(EVar "_14"%string);(EVar "_13"%string);(EVar "_12"%string);(EVar "_11"%string);(EVar "_10"%string)])]))]) |};
          {| identifier := ("rkeymerge3_1"%string, 10) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string;"_6"%string;"_7"%string;"_8"%string;"_9"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string);(EVar "_6"%string);(EVar "_7"%string);(EVar "_8"%string);(EVar "_9"%string)]) [([(PVar "I"%string);(PCons (PVar "H1"%string) (PVar "T1"%string));(PVar "M"%string);(PVar "D"%string);(PVar "E2"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "E3"%string);(PVar "H3"%string);(PVar "T3"%string)], (ELit (Atom "true"%string)), (ECase (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "I"%string);(EVar "H1"%string)]) [([(PVar "E1"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "E1"%string);(EVar "E2"%string)]), (ECase (EValues [(EVar "I"%string);(EVar "E1"%string);(EVar "H1"%string);(EVar "T1"%string);(EVar "E2"%string);(EVar "H2"%string);(EVar "T2"%string);(EVar "E3"%string);(EVar "H3"%string);(EVar "T3"%string);(EVar "M"%string);(EVar "T2"%string)]) [([(PVar "_34"%string);(PVar "_35"%string);(PVar "_36"%string);(PVar "_37"%string);(PVar "_38"%string);(PVar "_39"%string);(PVar "_40"%string);(PVar "_41"%string);(PVar "_42"%string);(PVar "_43"%string);(PVar "_44"%string);(PVar "_D"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "_38"%string);(EVar "_41"%string)]), (EApp (EFunId ("rkeymerge3_12_3"%string, 9)) [(EVar "_34"%string);(EVar "_35"%string);(EVar "_36"%string);(EVar "_37"%string);(EVar "_38"%string);(EVar "_39"%string);(EVar "_40"%string);(EVar "_43"%string);(ECons (EVar "_42"%string) (EVar "_44"%string))]));([(PVar "_45"%string);(PVar "_46"%string);(PVar "_47"%string);(PVar "_48"%string);(PVar "_E2"%string);(PVar "_49"%string);(PVar "_50"%string);(PVar "_51"%string);(PVar "_52"%string);(PVar "_53"%string);(PVar "_54"%string);(PVar "_55"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rkeymerge3_2"%string, 10)) [(EVar "_45"%string);(EVar "_46"%string);(EVar "_47"%string);(EVar "_48"%string);(EVar "_50"%string);(ECons (EVar "_49"%string) (EVar "_54"%string));(EVar "_55"%string);(EVar "_51"%string);(EVar "_52"%string);(EVar "_53"%string)]))]));([(PVar "E1"%string)], (ELit (Atom "true"%string)), (ECase (EValues [(EVar "I"%string);(EVar "E1"%string);(EVar "H1"%string);(EVar "T1"%string);(EVar "E2"%string);(EVar "H2"%string);(EVar "T2"%string);(EVar "E3"%string);(EVar "H3"%string);(EVar "T3"%string);(EVar "M"%string);(EVar "D"%string)]) [([(PVar "_66"%string);(PVar "_67"%string);(PVar "_68"%string);(PVar "_69"%string);(PVar "_70"%string);(PVar "_71"%string);(PVar "_72"%string);(PVar "_73"%string);(PVar "_74"%string);(PVar "_75"%string);(PVar "_76"%string);(PVar "_D"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "_67"%string);(EVar "_73"%string)]), (EApp (EFunId ("rkeymerge3_21_3"%string, 9)) [(EVar "_66"%string);(EVar "_67"%string);(EVar "_68"%string);(EVar "_69"%string);(EVar "_70"%string);(EVar "_71"%string);(EVar "_72"%string);(EVar "_75"%string);(ECons (EVar "_74"%string) (EVar "_76"%string))]));([(PVar "_77"%string);(PVar "_E1"%string);(PVar "_78"%string);(PVar "_79"%string);(PVar "_80"%string);(PVar "_81"%string);(PVar "_82"%string);(PVar "_83"%string);(PVar "_84"%string);(PVar "_85"%string);(PVar "_86"%string);(PVar "_87"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rkeymerge3_1"%string, 10)) [(EVar "_77"%string);(EVar "_79"%string);(ECons (EVar "_78"%string) (EVar "_86"%string));(EVar "_87"%string);(EVar "_80"%string);(EVar "_81"%string);(EVar "_82"%string);(EVar "_83"%string);(EVar "_84"%string);(EVar "_85"%string)]))]))]));([(PVar "I"%string);PNil;(PVar "M"%string);(PVar "_D"%string);(PVar "E2"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "E3"%string);(PVar "H3"%string);(PVar "T3"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "E2"%string);(EVar "E3"%string)]), (EApp (EFunId ("rkeymerge2_2"%string, 7)) [(EVar "I"%string);(EVar "E2"%string);(EVar "T2"%string);(EVar "H3"%string);(EVar "T3"%string);(EVar "M"%string);(EVar "H2"%string)]));([(PVar "I"%string);PNil;(PVar "M"%string);(PVar "_D"%string);(PVar "_E2"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "E3"%string);(PVar "H3"%string);(PVar "T3"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rkeymerge2_1"%string, 6)) [(EVar "I"%string);(EVar "T2"%string);(EVar "E3"%string);(EVar "H3"%string);(EVar "T3"%string);(ECons (EVar "H2"%string) (EVar "M"%string))]));([(PVar "_20"%string);(PVar "_19"%string);(PVar "_18"%string);(PVar "_17"%string);(PVar "_16"%string);(PVar "_15"%string);(PVar "_14"%string);(PVar "_13"%string);(PVar "_12"%string);(PVar "_11"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_20"%string);(EVar "_19"%string);(EVar "_18"%string);(EVar "_17"%string);(EVar "_16"%string);(EVar "_15"%string);(EVar "_14"%string);(EVar "_13"%string);(EVar "_12"%string);(EVar "_11"%string)])]))]) |};
          {| identifier := ("rkeymerge3_2"%string, 10) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string;"_6"%string;"_7"%string;"_8"%string;"_9"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string);(EVar "_6"%string);(EVar "_7"%string);(EVar "_8"%string);(EVar "_9"%string)]) [([(PVar "I"%string);(PVar "E1"%string);(PVar "H1"%string);(PVar "T1"%string);(PCons (PVar "H2"%string) (PVar "T2"%string));(PVar "M"%string);(PVar "D"%string);(PVar "E3"%string);(PVar "H3"%string);(PVar "T3"%string)], (ELit (Atom "true"%string)), (ECase (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "I"%string);(EVar "H2"%string)]) [([(PVar "E2"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "E1"%string);(EVar "E2"%string)]), (ECase (EValues [(EVar "I"%string);(EVar "E1"%string);(EVar "H1"%string);(EVar "T1"%string);(EVar "E2"%string);(EVar "H2"%string);(EVar "T2"%string);(EVar "E3"%string);(EVar "H3"%string);(EVar "T3"%string);(EVar "M"%string);(EVar "D"%string)]) [([(PVar "_34"%string);(PVar "_35"%string);(PVar "_36"%string);(PVar "_37"%string);(PVar "_38"%string);(PVar "_39"%string);(PVar "_40"%string);(PVar "_41"%string);(PVar "_42"%string);(PVar "_43"%string);(PVar "_44"%string);(PVar "_D"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "_38"%string);(EVar "_41"%string)]), (EApp (EFunId ("rkeymerge3_12_3"%string, 9)) [(EVar "_34"%string);(EVar "_35"%string);(EVar "_36"%string);(EVar "_37"%string);(EVar "_38"%string);(EVar "_39"%string);(EVar "_40"%string);(EVar "_43"%string);(ECons (EVar "_42"%string) (EVar "_44"%string))]));([(PVar "_45"%string);(PVar "_46"%string);(PVar "_47"%string);(PVar "_48"%string);(PVar "_E2"%string);(PVar "_49"%string);(PVar "_50"%string);(PVar "_51"%string);(PVar "_52"%string);(PVar "_53"%string);(PVar "_54"%string);(PVar "_55"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rkeymerge3_2"%string, 10)) [(EVar "_45"%string);(EVar "_46"%string);(EVar "_47"%string);(EVar "_48"%string);(EVar "_50"%string);(ECons (EVar "_49"%string) (EVar "_54"%string));(EVar "_55"%string);(EVar "_51"%string);(EVar "_52"%string);(EVar "_53"%string)]))]));([(PVar "E2"%string)], (ELit (Atom "true"%string)), (ECase (EValues [(EVar "I"%string);(EVar "E1"%string);(EVar "H1"%string);(EVar "T1"%string);(EVar "E2"%string);(EVar "H2"%string);(EVar "T2"%string);(EVar "E3"%string);(EVar "H3"%string);(EVar "T3"%string);(EVar "M"%string);(EVar "T1"%string)]) [([(PVar "_66"%string);(PVar "_67"%string);(PVar "_68"%string);(PVar "_69"%string);(PVar "_70"%string);(PVar "_71"%string);(PVar "_72"%string);(PVar "_73"%string);(PVar "_74"%string);(PVar "_75"%string);(PVar "_76"%string);(PVar "_D"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "_67"%string);(EVar "_73"%string)]), (EApp (EFunId ("rkeymerge3_21_3"%string, 9)) [(EVar "_66"%string);(EVar "_67"%string);(EVar "_68"%string);(EVar "_69"%string);(EVar "_70"%string);(EVar "_71"%string);(EVar "_72"%string);(EVar "_75"%string);(ECons (EVar "_74"%string) (EVar "_76"%string))]));([(PVar "_77"%string);(PVar "_E1"%string);(PVar "_78"%string);(PVar "_79"%string);(PVar "_80"%string);(PVar "_81"%string);(PVar "_82"%string);(PVar "_83"%string);(PVar "_84"%string);(PVar "_85"%string);(PVar "_86"%string);(PVar "_87"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rkeymerge3_1"%string, 10)) [(EVar "_77"%string);(EVar "_79"%string);(ECons (EVar "_78"%string) (EVar "_86"%string));(EVar "_87"%string);(EVar "_80"%string);(EVar "_81"%string);(EVar "_82"%string);(EVar "_83"%string);(EVar "_84"%string);(EVar "_85"%string)]))]))]));([(PVar "I"%string);(PVar "E1"%string);(PVar "H1"%string);(PVar "T1"%string);PNil;(PVar "M"%string);(PVar "_D"%string);(PVar "E3"%string);(PVar "H3"%string);(PVar "T3"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "E1"%string);(EVar "E3"%string)]), (EApp (EFunId ("rkeymerge2_2"%string, 7)) [(EVar "I"%string);(EVar "E1"%string);(EVar "T1"%string);(EVar "H3"%string);(EVar "T3"%string);(EVar "M"%string);(EVar "H1"%string)]));([(PVar "I"%string);(PVar "_E1"%string);(PVar "H1"%string);(PVar "T1"%string);PNil;(PVar "M"%string);(PVar "_D"%string);(PVar "E3"%string);(PVar "H3"%string);(PVar "T3"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rkeymerge2_1"%string, 6)) [(EVar "I"%string);(EVar "T1"%string);(EVar "E3"%string);(EVar "H3"%string);(EVar "T3"%string);(ECons (EVar "H1"%string) (EVar "M"%string))]));([(PVar "_20"%string);(PVar "_19"%string);(PVar "_18"%string);(PVar "_17"%string);(PVar "_16"%string);(PVar "_15"%string);(PVar "_14"%string);(PVar "_13"%string);(PVar "_12"%string);(PVar "_11"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_20"%string);(EVar "_19"%string);(EVar "_18"%string);(EVar "_17"%string);(EVar "_16"%string);(EVar "_15"%string);(EVar "_14"%string);(EVar "_13"%string);(EVar "_12"%string);(EVar "_11"%string)])]))]) |};
          {| identifier := ("rkeymerge3_12"%string, 12) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string;"_6"%string;"_7"%string;"_8"%string;"_9"%string;"_10"%string;"_11"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string);(EVar "_6"%string);(EVar "_7"%string);(EVar "_8"%string);(EVar "_9"%string);(EVar "_10"%string);(EVar "_11"%string)]) [([(PVar "I"%string);(PVar "E1"%string);(PVar "H1"%string);(PVar "T1"%string);(PVar "E2"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "E3"%string);(PVar "H3"%string);(PVar "T3"%string);(PVar "M"%string);(PVar "_D"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "E2"%string);(EVar "E3"%string)]), (EApp (EFunId ("rkeymerge3_12_3"%string, 9)) [(EVar "I"%string);(EVar "E1"%string);(EVar "H1"%string);(EVar "T1"%string);(EVar "E2"%string);(EVar "H2"%string);(EVar "T2"%string);(EVar "T3"%string);(ECons (EVar "H3"%string) (EVar "M"%string))]));([(PVar "I"%string);(PVar "E1"%string);(PVar "H1"%string);(PVar "T1"%string);(PVar "_E2"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "E3"%string);(PVar "H3"%string);(PVar "T3"%string);(PVar "M"%string);(PVar "D"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rkeymerge3_2"%string, 10)) [(EVar "I"%string);(EVar "E1"%string);(EVar "H1"%string);(EVar "T1"%string);(EVar "T2"%string);(ECons (EVar "H2"%string) (EVar "M"%string));(EVar "D"%string);(EVar "E3"%string);(EVar "H3"%string);(EVar "T3"%string)]))]) |};
          {| identifier := ("rkeymerge3_12_3"%string, 9) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string;"_6"%string;"_7"%string;"_8"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string);(EVar "_6"%string);(EVar "_7"%string);(EVar "_8"%string)]) [([(PVar "I"%string);(PVar "E1"%string);(PVar "H1"%string);(PVar "T1"%string);(PVar "E2"%string);(PVar "H2"%string);(PVar "T2"%string);(PCons (PVar "H3"%string) (PVar "T3"%string));(PVar "M"%string)], (ELit (Atom "true"%string)), (ECase (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "I"%string);(EVar "H3"%string)]) [([(PVar "E3"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "E2"%string);(EVar "E3"%string)]), (EApp (EFunId ("rkeymerge3_12_3"%string, 9)) [(EVar "I"%string);(EVar "E1"%string);(EVar "H1"%string);(EVar "T1"%string);(EVar "E2"%string);(EVar "H2"%string);(EVar "T2"%string);(EVar "T3"%string);(ECons (EVar "H3"%string) (EVar "M"%string))]));([(PVar "E3"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rkeymerge3_2"%string, 10)) [(EVar "I"%string);(EVar "E1"%string);(EVar "H1"%string);(EVar "T1"%string);(EVar "T2"%string);(ECons (EVar "H2"%string) (EVar "M"%string));(EVar "T2"%string);(EVar "E3"%string);(EVar "H3"%string);(EVar "T3"%string)]))]));([(PVar "I"%string);(PVar "E1"%string);(PVar "H1"%string);(PVar "T1"%string);(PVar "_E2"%string);(PVar "H2"%string);(PVar "T2"%string);PNil;(PVar "M"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rkeymerge2_2"%string, 7)) [(EVar "I"%string);(EVar "E1"%string);(EVar "T1"%string);(EVar "H2"%string);(EVar "T2"%string);(EVar "M"%string);(EVar "H1"%string)]));([(PVar "_18"%string);(PVar "_17"%string);(PVar "_16"%string);(PVar "_15"%string);(PVar "_14"%string);(PVar "_13"%string);(PVar "_12"%string);(PVar "_11"%string);(PVar "_10"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_18"%string);(EVar "_17"%string);(EVar "_16"%string);(EVar "_15"%string);(EVar "_14"%string);(EVar "_13"%string);(EVar "_12"%string);(EVar "_11"%string);(EVar "_10"%string)])]))]) |};
          {| identifier := ("rkeymerge3_21"%string, 12) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string;"_6"%string;"_7"%string;"_8"%string;"_9"%string;"_10"%string;"_11"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string);(EVar "_6"%string);(EVar "_7"%string);(EVar "_8"%string);(EVar "_9"%string);(EVar "_10"%string);(EVar "_11"%string)]) [([(PVar "I"%string);(PVar "E1"%string);(PVar "H1"%string);(PVar "T1"%string);(PVar "E2"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "E3"%string);(PVar "H3"%string);(PVar "T3"%string);(PVar "M"%string);(PVar "_D"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "E1"%string);(EVar "E3"%string)]), (EApp (EFunId ("rkeymerge3_21_3"%string, 9)) [(EVar "I"%string);(EVar "E1"%string);(EVar "H1"%string);(EVar "T1"%string);(EVar "E2"%string);(EVar "H2"%string);(EVar "T2"%string);(EVar "T3"%string);(ECons (EVar "H3"%string) (EVar "M"%string))]));([(PVar "I"%string);(PVar "_E1"%string);(PVar "H1"%string);(PVar "T1"%string);(PVar "E2"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "E3"%string);(PVar "H3"%string);(PVar "T3"%string);(PVar "M"%string);(PVar "D"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rkeymerge3_1"%string, 10)) [(EVar "I"%string);(EVar "T1"%string);(ECons (EVar "H1"%string) (EVar "M"%string));(EVar "D"%string);(EVar "E2"%string);(EVar "H2"%string);(EVar "T2"%string);(EVar "E3"%string);(EVar "H3"%string);(EVar "T3"%string)]))]) |};
          {| identifier := ("rkeymerge3_21_3"%string, 9) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string;"_6"%string;"_7"%string;"_8"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string);(EVar "_6"%string);(EVar "_7"%string);(EVar "_8"%string)]) [([(PVar "I"%string);(PVar "E1"%string);(PVar "H1"%string);(PVar "T1"%string);(PVar "E2"%string);(PVar "H2"%string);(PVar "T2"%string);(PCons (PVar "H3"%string) (PVar "T3"%string));(PVar "M"%string)], (ELit (Atom "true"%string)), (ECase (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "I"%string);(EVar "H3"%string)]) [([(PVar "E3"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "E1"%string);(EVar "E3"%string)]), (EApp (EFunId ("rkeymerge3_21_3"%string, 9)) [(EVar "I"%string);(EVar "E1"%string);(EVar "H1"%string);(EVar "T1"%string);(EVar "E2"%string);(EVar "H2"%string);(EVar "T2"%string);(EVar "T3"%string);(ECons (EVar "H3"%string) (EVar "M"%string))]));([(PVar "E3"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rkeymerge3_1"%string, 10)) [(EVar "I"%string);(EVar "T1"%string);(ECons (EVar "H1"%string) (EVar "M"%string));(EVar "T1"%string);(EVar "E2"%string);(EVar "H2"%string);(EVar "T2"%string);(EVar "E3"%string);(EVar "H3"%string);(EVar "T3"%string)]))]));([(PVar "I"%string);(PVar "_E1"%string);(PVar "H1"%string);(PVar "T1"%string);(PVar "E2"%string);(PVar "H2"%string);(PVar "T2"%string);PNil;(PVar "M"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rkeymerge2_1"%string, 6)) [(EVar "I"%string);(EVar "T1"%string);(EVar "E2"%string);(EVar "H2"%string);(EVar "T2"%string);(ECons (EVar "H1"%string) (EVar "M"%string))]));([(PVar "_18"%string);(PVar "_17"%string);(PVar "_16"%string);(PVar "_15"%string);(PVar "_14"%string);(PVar "_13"%string);(PVar "_12"%string);(PVar "_11"%string);(PVar "_10"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_18"%string);(EVar "_17"%string);(EVar "_16"%string);(EVar "_15"%string);(EVar "_14"%string);(EVar "_13"%string);(EVar "_12"%string);(EVar "_11"%string);(EVar "_10"%string)])]))]) |};
          {| identifier := ("keymerge2_1"%string, 6) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string)]) [([(PVar "I"%string);(PCons (PVar "H1"%string) (PVar "T1"%string));(PVar "E2"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "M"%string)], (ELit (Atom "true"%string)), (ECase (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "I"%string);(EVar "H1"%string)]) [([(PVar "E1"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "E1"%string);(EVar "E2"%string)]), (EApp (EFunId ("keymerge2_1"%string, 6)) [(EVar "I"%string);(EVar "T1"%string);(EVar "E2"%string);(EVar "H2"%string);(EVar "T2"%string);(ECons (EVar "H1"%string) (EVar "M"%string))]));([(PVar "E1"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("keymerge2_2"%string, 7)) [(EVar "I"%string);(EVar "T1"%string);(EVar "E1"%string);(EVar "H2"%string);(EVar "T2"%string);(EVar "M"%string);(EVar "H1"%string)]))]));([(PVar "_I"%string);PNil;(PVar "_E2"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "M"%string)], (ELit (Atom "true"%string)), (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "T2"%string);(ECons (EVar "H2"%string) (EVar "M"%string))]));([(PVar "_12"%string);(PVar "_11"%string);(PVar "_10"%string);(PVar "_9"%string);(PVar "_8"%string);(PVar "_7"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_12"%string);(EVar "_11"%string);(EVar "_10"%string);(EVar "_9"%string);(EVar "_8"%string);(EVar "_7"%string)])]))]) |};
          {| identifier := ("keymerge2_2"%string, 7) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string;"_6"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string);(EVar "_6"%string)]) [([(PVar "I"%string);(PVar "T1"%string);(PVar "E1"%string);(PVar "HdM"%string);(PCons (PVar "H2"%string) (PVar "T2"%string));(PVar "M"%string);(PVar "H1"%string)], (ELit (Atom "true"%string)), (ECase (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "I"%string);(EVar "H2"%string)]) [([(PVar "E2"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "E1"%string);(EVar "E2"%string)]), (EApp (EFunId ("keymerge2_1"%string, 6)) [(EVar "I"%string);(EVar "T1"%string);(EVar "E2"%string);(EVar "H2"%string);(EVar "T2"%string);(ECons (EVar "H1"%string) (ECons (EVar "HdM"%string) (EVar "M"%string)))]));([(PVar "_E2"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("keymerge2_2"%string, 7)) [(EVar "I"%string);(EVar "T1"%string);(EVar "E1"%string);(EVar "H2"%string);(EVar "T2"%string);(ECons (EVar "HdM"%string) (EVar "M"%string));(EVar "H1"%string)]))]));([(PVar "_I"%string);(PVar "T1"%string);(PVar "_E1"%string);(PVar "HdM"%string);PNil;(PVar "M"%string);(PVar "H1"%string)], (ELit (Atom "true"%string)), (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "T1"%string);(ECons (EVar "H1"%string) (ECons (EVar "HdM"%string) (EVar "M"%string)))]));([(PVar "_14"%string);(PVar "_13"%string);(PVar "_12"%string);(PVar "_11"%string);(PVar "_10"%string);(PVar "_9"%string);(PVar "_8"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_14"%string);(EVar "_13"%string);(EVar "_12"%string);(EVar "_11"%string);(EVar "_10"%string);(EVar "_9"%string);(EVar "_8"%string)])]))]) |};
          {| identifier := ("rkeymerge2_1"%string, 6) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string)]) [([(PVar "I"%string);(PCons (PVar "H1"%string) (PVar "T1"%string));(PVar "E2"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "M"%string)], (ELit (Atom "true"%string)), (ECase (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "I"%string);(EVar "H1"%string)]) [([(PVar "E1"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "E1"%string);(EVar "E2"%string)]), (EApp (EFunId ("rkeymerge2_2"%string, 7)) [(EVar "I"%string);(EVar "E1"%string);(EVar "T1"%string);(EVar "H2"%string);(EVar "T2"%string);(EVar "M"%string);(EVar "H1"%string)]));([(PVar "_E1"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rkeymerge2_1"%string, 6)) [(EVar "I"%string);(EVar "T1"%string);(EVar "E2"%string);(EVar "H2"%string);(EVar "T2"%string);(ECons (EVar "H1"%string) (EVar "M"%string))]))]));([(PVar "_I"%string);PNil;(PVar "_E2"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "M"%string)], (ELit (Atom "true"%string)), (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "T2"%string);(ECons (EVar "H2"%string) (EVar "M"%string))]));([(PVar "_12"%string);(PVar "_11"%string);(PVar "_10"%string);(PVar "_9"%string);(PVar "_8"%string);(PVar "_7"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_12"%string);(EVar "_11"%string);(EVar "_10"%string);(EVar "_9"%string);(EVar "_8"%string);(EVar "_7"%string)])]))]) |};
          {| identifier := ("rkeymerge2_2"%string, 7) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string;"_6"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string);(EVar "_6"%string)]) [([(PVar "I"%string);(PVar "E1"%string);(PVar "T1"%string);(PVar "HdM"%string);(PCons (PVar "H2"%string) (PVar "T2"%string));(PVar "M"%string);(PVar "H1"%string)], (ELit (Atom "true"%string)), (ECase (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "I"%string);(EVar "H2"%string)]) [([(PVar "E2"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "E1"%string);(EVar "E2"%string)]), (EApp (EFunId ("rkeymerge2_2"%string, 7)) [(EVar "I"%string);(EVar "E1"%string);(EVar "T1"%string);(EVar "H2"%string);(EVar "T2"%string);(ECons (EVar "HdM"%string) (EVar "M"%string));(EVar "H1"%string)]));([(PVar "E2"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rkeymerge2_1"%string, 6)) [(EVar "I"%string);(EVar "T1"%string);(EVar "E2"%string);(EVar "H2"%string);(EVar "T2"%string);(ECons (EVar "H1"%string) (ECons (EVar "HdM"%string) (EVar "M"%string)))]))]));([(PVar "_I"%string);(PVar "_E1"%string);(PVar "T1"%string);(PVar "HdM"%string);PNil;(PVar "M"%string);(PVar "H1"%string)], (ELit (Atom "true"%string)), (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "T1"%string);(ECons (EVar "H1"%string) (ECons (EVar "HdM"%string) (EVar "M"%string)))]));([(PVar "_14"%string);(PVar "_13"%string);(PVar "_12"%string);(PVar "_11"%string);(PVar "_10"%string);(PVar "_9"%string);(PVar "_8"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_14"%string);(EVar "_13"%string);(EVar "_12"%string);(EVar "_11"%string);(EVar "_10"%string);(EVar "_9"%string);(EVar "_8"%string)])]))]) |};
          {| identifier := ("ukeysplit_1"%string, 8) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string;"_6"%string;"_7"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string);(EVar "_6"%string);(EVar "_7"%string)]) [([(PVar "I"%string);(PVar "X"%string);(PVar "EX"%string);(PVar "Y"%string);(PVar "EY"%string);(PCons (PVar "Z"%string) (PVar "L"%string));(PVar "R"%string);(PVar "Rs"%string)], (ELit (Atom "true"%string)), (ECase (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "I"%string);(EVar "Z"%string)]) [([(PVar "EZ"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "EY"%string);(EVar "EZ"%string)]), (EApp (EFunId ("ukeysplit_1"%string, 8)) [(EVar "I"%string);(EVar "X"%string);(EVar "EX"%string);(EVar "Y"%string);(EVar "EY"%string);(EVar "L"%string);(EVar "R"%string);(EVar "Rs"%string)]));([(PVar "EZ"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "<"%string)) [(EVar "EY"%string);(EVar "EZ"%string)]), (EApp (EFunId ("ukeysplit_1"%string, 8)) [(EVar "I"%string);(EVar "Y"%string);(EVar "EY"%string);(EVar "Z"%string);(EVar "EZ"%string);(EVar "L"%string);(ECons (EVar "X"%string) (EVar "R"%string));(EVar "Rs"%string)]));([(PVar "EZ"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "EX"%string);(EVar "EZ"%string)]), (EApp (EFunId ("ukeysplit_1"%string, 8)) [(EVar "I"%string);(EVar "X"%string);(EVar "EX"%string);(EVar "Y"%string);(EVar "EY"%string);(EVar "L"%string);(EVar "R"%string);(EVar "Rs"%string)]));([(PVar "EZ"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "<"%string)) [(EVar "EX"%string);(EVar "EZ"%string)]), (EApp (EFunId ("ukeysplit_1"%string, 8)) [(EVar "I"%string);(EVar "Z"%string);(EVar "EZ"%string);(EVar "Y"%string);(EVar "EY"%string);(EVar "L"%string);(ECons (EVar "X"%string) (EVar "R"%string));(EVar "Rs"%string)]));([(PVar "_EZ"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "R"%string);ENil]), (EApp (EFunId ("ukeysplit_1"%string, 8)) [(EVar "I"%string);(EVar "X"%string);(EVar "EX"%string);(EVar "Y"%string);(EVar "EY"%string);(EVar "L"%string);(ECons (EVar "Z"%string) ENil);(EVar "Rs"%string)]));([(PVar "EZ"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("ukeysplit_1_1"%string, 10)) [(EVar "I"%string);(EVar "X"%string);(EVar "EX"%string);(EVar "Y"%string);(EVar "EY"%string);(EVar "L"%string);(EVar "R"%string);(EVar "Rs"%string);(EVar "Z"%string);(EVar "EZ"%string)]))]));([(PVar "I"%string);(PVar "X"%string);(PVar "_EX"%string);(PVar "Y"%string);(PVar "_EY"%string);PNil;(PVar "R"%string);(PVar "Rs"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rukeymergel"%string, 3)) [(EVar "I"%string);(ECons (ECons (EVar "Y"%string) (ECons (EVar "X"%string) (EVar "R"%string))) (EVar "Rs"%string));ENil]));([(PVar "_16"%string);(PVar "_15"%string);(PVar "_14"%string);(PVar "_13"%string);(PVar "_12"%string);(PVar "_11"%string);(PVar "_10"%string);(PVar "_9"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_16"%string);(EVar "_15"%string);(EVar "_14"%string);(EVar "_13"%string);(EVar "_12"%string);(EVar "_11"%string);(EVar "_10"%string);(EVar "_9"%string)])]))]) |};
          {| identifier := ("ukeysplit_1_1"%string, 10) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string;"_6"%string;"_7"%string;"_8"%string;"_9"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string);(EVar "_6"%string);(EVar "_7"%string);(EVar "_8"%string);(EVar "_9"%string)]) [([(PVar "I"%string);(PVar "X"%string);(PVar "EX"%string);(PVar "Y"%string);(PVar "EY"%string);(PCons (PVar "Z"%string) (PVar "L"%string));(PVar "R"%string);(PVar "Rs"%string);(PVar "S"%string);(PVar "ES"%string)], (ELit (Atom "true"%string)), (ECase (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "I"%string);(EVar "Z"%string)]) [([(PVar "EZ"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "EY"%string);(EVar "EZ"%string)]), (EApp (EFunId ("ukeysplit_1_1"%string, 10)) [(EVar "I"%string);(EVar "X"%string);(EVar "EX"%string);(EVar "Y"%string);(EVar "EY"%string);(EVar "L"%string);(EVar "R"%string);(EVar "Rs"%string);(EVar "S"%string);(EVar "ES"%string)]));([(PVar "EZ"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "<"%string)) [(EVar "EY"%string);(EVar "EZ"%string)]), (EApp (EFunId ("ukeysplit_1_1"%string, 10)) [(EVar "I"%string);(EVar "Y"%string);(EVar "EY"%string);(EVar "Z"%string);(EVar "EZ"%string);(EVar "L"%string);(ECons (EVar "X"%string) (EVar "R"%string));(EVar "Rs"%string);(EVar "S"%string);(EVar "ES"%string)]));([(PVar "EZ"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "EX"%string);(EVar "EZ"%string)]), (EApp (EFunId ("ukeysplit_1_1"%string, 10)) [(EVar "I"%string);(EVar "X"%string);(EVar "EX"%string);(EVar "Y"%string);(EVar "EY"%string);(EVar "L"%string);(EVar "R"%string);(EVar "Rs"%string);(EVar "S"%string);(EVar "ES"%string)]));([(PVar "EZ"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "<"%string)) [(EVar "EX"%string);(EVar "EZ"%string)]), (EApp (EFunId ("ukeysplit_1_1"%string, 10)) [(EVar "I"%string);(EVar "Z"%string);(EVar "EZ"%string);(EVar "Y"%string);(EVar "EY"%string);(EVar "L"%string);(ECons (EVar "X"%string) (EVar "R"%string));(EVar "Rs"%string);(EVar "S"%string);(EVar "ES"%string)]));([(PVar "EZ"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "ES"%string);(EVar "EZ"%string)]), (EApp (EFunId ("ukeysplit_1_1"%string, 10)) [(EVar "I"%string);(EVar "X"%string);(EVar "EX"%string);(EVar "Y"%string);(EVar "EY"%string);(EVar "L"%string);(EVar "R"%string);(EVar "Rs"%string);(EVar "S"%string);(EVar "ES"%string)]));([(PVar "EZ"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "<"%string)) [(EVar "ES"%string);(EVar "EZ"%string)]), (EApp (EFunId ("ukeysplit_1"%string, 8)) [(EVar "I"%string);(EVar "S"%string);(EVar "ES"%string);(EVar "Z"%string);(EVar "EZ"%string);(EVar "L"%string);ENil;(ECons (ECons (EVar "Y"%string) (ECons (EVar "X"%string) (EVar "R"%string))) (EVar "Rs"%string))]));([(PVar "EZ"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("ukeysplit_1"%string, 8)) [(EVar "I"%string);(EVar "Z"%string);(EVar "EZ"%string);(EVar "S"%string);(EVar "ES"%string);(EVar "L"%string);ENil;(ECons (ECons (EVar "Y"%string) (ECons (EVar "X"%string) (EVar "R"%string))) (EVar "Rs"%string))]))]));([(PVar "I"%string);(PVar "X"%string);(PVar "_EX"%string);(PVar "Y"%string);(PVar "_EY"%string);PNil;(PVar "R"%string);(PVar "Rs"%string);(PVar "S"%string);(PVar "_ES"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rukeymergel"%string, 3)) [(EVar "I"%string);(ECons (ECons (EVar "S"%string) ENil) (ECons (ECons (EVar "Y"%string) (ECons (EVar "X"%string) (EVar "R"%string))) (EVar "Rs"%string)));ENil]));([(PVar "_20"%string);(PVar "_19"%string);(PVar "_18"%string);(PVar "_17"%string);(PVar "_16"%string);(PVar "_15"%string);(PVar "_14"%string);(PVar "_13"%string);(PVar "_12"%string);(PVar "_11"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_20"%string);(EVar "_19"%string);(EVar "_18"%string);(EVar "_17"%string);(EVar "_16"%string);(EVar "_15"%string);(EVar "_14"%string);(EVar "_13"%string);(EVar "_12"%string);(EVar "_11"%string)])]))]) |};
          {| identifier := ("ukeysplit_2"%string, 5) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string)]) [([(PVar "I"%string);(PVar "Y"%string);(PVar "EY"%string);(PCons (PVar "Z"%string) (PVar "L"%string));(PVar "R"%string)], (ELit (Atom "true"%string)), (ECase (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "I"%string);(EVar "Z"%string)]) [([(PVar "EZ"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "EY"%string);(EVar "EZ"%string)]), (EApp (EFunId ("ukeysplit_2"%string, 5)) [(EVar "I"%string);(EVar "Y"%string);(EVar "EY"%string);(EVar "L"%string);(EVar "R"%string)]));([(PVar "EZ"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "<"%string)) [(EVar "EY"%string);(EVar "EZ"%string)]), (ELet ["_5"%string] (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "R"%string);ENil]) (EApp (EFunId ("ukeysplit_1"%string, 8)) [(EVar "I"%string);(EVar "Y"%string);(EVar "EY"%string);(EVar "Z"%string);(EVar "EZ"%string);(EVar "L"%string);ENil;(ECons (EVar "_5"%string) ENil)])));([(PVar "EZ"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("ukeysplit_2"%string, 5)) [(EVar "I"%string);(EVar "Z"%string);(EVar "EZ"%string);(EVar "L"%string);(ECons (EVar "Y"%string) (EVar "R"%string))]))]));([(PVar "_I"%string);(PVar "Y"%string);(PVar "_EY"%string);PNil;(PVar "R"%string)], (ELit (Atom "true"%string)), (ECons (EVar "Y"%string) (EVar "R"%string)));([(PVar "_11"%string);(PVar "_10"%string);(PVar "_9"%string);(PVar "_8"%string);(PVar "_7"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_11"%string);(EVar "_10"%string);(EVar "_9"%string);(EVar "_8"%string);(EVar "_7"%string)])]))]) |};
          {| identifier := ("ukeymergel"%string, 3) ; varl := ["_0"%string;"_1"%string;"_2"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string)]) [([(PVar "I"%string);(PCons (PVar "T1"%string) (PCons (PCons (PVar "H2"%string) (PVar "T2"%string)) (PCons (PCons (PVar "H3"%string) (PVar "T3"%string)) (PVar "L"%string))));(PVar "Acc"%string)], (ELit (Atom "true"%string)), (ELet ["_4"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "I"%string);(EVar "H2"%string)]) (ELet ["_3"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "I"%string);(EVar "H3"%string)]) (ELet ["M"%string] (EApp (EFunId ("ukeymerge3_1"%string, 11)) [(EVar "I"%string);(EVar "T1"%string);(EVar "Acc"%string);(ECons (EVar "H2"%string) (EVar "H3"%string));(EVar "_4"%string);(EVar "H2"%string);(EVar "T2"%string);ENil;(EVar "_3"%string);(EVar "H3"%string);(EVar "T3"%string)]) (EApp (EFunId ("ukeymergel"%string, 3)) [(EVar "I"%string);(EVar "L"%string);(ECons (EVar "M"%string) (EVar "Acc"%string))])))));([(PVar "I"%string);(PCons (PCons (PVar "H1"%string) (PVar "T1"%string)) (PCons (PVar "T2"%string) (PVar "L"%string)));(PVar "Acc"%string)], (ELit (Atom "true"%string)), (ELet ["_6"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "I"%string);(EVar "H1"%string)]) (ELet ["_7"%string] (EApp (EFunId ("ukeymerge2_2"%string, 6)) [(EVar "I"%string);(EVar "T1"%string);(EVar "_6"%string);(EVar "H1"%string);(EVar "T2"%string);ENil]) (EApp (EFunId ("ukeymergel"%string, 3)) [(EVar "I"%string);(EVar "L"%string);(ECons (EVar "_7"%string) (EVar "Acc"%string))]))));([(PVar "_I"%string);(PCons (PVar "L"%string) PNil);PNil], (ELit (Atom "true"%string)), (EVar "L"%string));([(PVar "I"%string);(PCons (PVar "L"%string) PNil);(PVar "Acc"%string)], (ELit (Atom "true"%string)), (ELet ["_8"%string] (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "L"%string);ENil]) (EApp (EFunId ("rukeymergel"%string, 3)) [(EVar "I"%string);(ECons (EVar "_8"%string) (EVar "Acc"%string));ENil])));([(PVar "I"%string);PNil;(PVar "Acc"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rukeymergel"%string, 3)) [(EVar "I"%string);(EVar "Acc"%string);ENil]));([(PVar "_11"%string);(PVar "_10"%string);(PVar "_9"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_11"%string);(EVar "_10"%string);(EVar "_9"%string)])]))]) |};
          {| identifier := ("rukeymergel"%string, 3) ; varl := ["_0"%string;"_1"%string;"_2"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string)]) [([(PVar "I"%string);(PCons (PCons (PVar "H3"%string) (PVar "T3"%string)) (PCons (PCons (PVar "H2"%string) (PVar "T2"%string)) (PCons (PVar "T1"%string) (PVar "L"%string))));(PVar "Acc"%string)], (ELit (Atom "true"%string)), (ELet ["_4"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "I"%string);(EVar "H2"%string)]) (ELet ["_3"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "I"%string);(EVar "H3"%string)]) (ELet ["M"%string] (EApp (EFunId ("rukeymerge3_1"%string, 11)) [(EVar "I"%string);(EVar "T1"%string);(EVar "Acc"%string);ENil;(EVar "_4"%string);(EVar "H2"%string);(EVar "T2"%string);ENil;(EVar "_3"%string);(EVar "H3"%string);(EVar "T3"%string)]) (EApp (EFunId ("rukeymergel"%string, 3)) [(EVar "I"%string);(EVar "L"%string);(ECons (EVar "M"%string) (EVar "Acc"%string))])))));([(PVar "I"%string);(PCons (PCons (PVar "H2"%string) (PVar "T2"%string)) (PCons (PVar "T1"%string) (PVar "L"%string)));(PVar "Acc"%string)], (ELit (Atom "true"%string)), (ELet ["_6"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "I"%string);(EVar "H2"%string)]) (ELet ["_7"%string] (EApp (EFunId ("rukeymerge2_1"%string, 6)) [(EVar "I"%string);(EVar "T1"%string);(EVar "_6"%string);(EVar "T2"%string);ENil;(EVar "H2"%string)]) (EApp (EFunId ("rukeymergel"%string, 3)) [(EVar "I"%string);(EVar "L"%string);(ECons (EVar "_7"%string) (EVar "Acc"%string))]))));([(PVar "I"%string);(PCons (PVar "L"%string) PNil);(PVar "Acc"%string)], (ELit (Atom "true"%string)), (ELet ["_8"%string] (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "L"%string);ENil]) (EApp (EFunId ("ukeymergel"%string, 3)) [(EVar "I"%string);(ECons (EVar "_8"%string) (EVar "Acc"%string));ENil])));([(PVar "I"%string);PNil;(PVar "Acc"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("ukeymergel"%string, 3)) [(EVar "I"%string);(EVar "Acc"%string);ENil]));([(PVar "_11"%string);(PVar "_10"%string);(PVar "_9"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_11"%string);(EVar "_10"%string);(EVar "_9"%string)])]))]) |};
          {| identifier := ("ukeymerge3_1"%string, 11) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string;"_6"%string;"_7"%string;"_8"%string;"_9"%string;"_10"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string);(EVar "_6"%string);(EVar "_7"%string);(EVar "_8"%string);(EVar "_9"%string);(EVar "_10"%string)]) [([(PVar "I"%string);(PCons (PVar "H1"%string) (PVar "T1"%string));(PVar "D"%string);(PVar "HdM"%string);(PVar "E2"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "M"%string);(PVar "E3"%string);(PVar "H3"%string);(PVar "T3"%string)], (ELit (Atom "true"%string)), (ECase (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "I"%string);(EVar "H1"%string)]) [([(PVar "E1"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "E1"%string);(EVar "E2"%string)]), (ECase (EValues [(EVar "I"%string);(EVar "E1"%string);(EVar "T1"%string);(EVar "H1"%string);(EVar "E2"%string);(EVar "H2"%string);(EVar "T2"%string);(EVar "E3"%string);(EVar "H3"%string);(EVar "T3"%string);(EVar "M"%string);(EVar "HdM"%string);(EVar "D"%string)]) [([(PVar "_37"%string);(PVar "_38"%string);(PVar "_39"%string);(PVar "_40"%string);(PVar "_41"%string);(PVar "_42"%string);(PVar "_43"%string);(PVar "_44"%string);(PVar "_45"%string);(PVar "_46"%string);(PVar "_47"%string);(PVar "_HdM"%string);(PVar "_48"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "_38"%string);(EVar "_44"%string)]), (EApp (EFunId ("ukeymerge3_1"%string, 11)) [(EVar "_37"%string);(EVar "_39"%string);(EVar "_48"%string);(EVar "_38"%string);(EVar "_41"%string);(EVar "_42"%string);(EVar "_43"%string);(ECons (EVar "_40"%string) (EVar "_47"%string));(EVar "_44"%string);(EVar "_45"%string);(EVar "_46"%string)]));([(PVar "_49"%string);(PVar "_50"%string);(PVar "_51"%string);(PVar "_52"%string);(PVar "_53"%string);(PVar "_54"%string);(PVar "_55"%string);(PVar "_56"%string);(PVar "_H3"%string);(PVar "_57"%string);(PVar "_58"%string);(PVar "_59"%string);(PVar "_D"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "_56"%string);(EVar "_59"%string)]), (EApp (EFunId ("ukeymerge3_12_3"%string, 9)) [(EVar "_49"%string);(EVar "_50"%string);(EVar "_51"%string);(EVar "_52"%string);(EVar "_53"%string);(EVar "_54"%string);(EVar "_55"%string);(EVar "_58"%string);(EVar "_57"%string)]));([(PVar "_60"%string);(PVar "_61"%string);(PVar "_62"%string);(PVar "_63"%string);(PVar "_64"%string);(PVar "_65"%string);(PVar "_66"%string);(PVar "_E3"%string);(PVar "_67"%string);(PVar "_68"%string);(PVar "_69"%string);(PVar "_HdM"%string);(PVar "_D"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("ukeymerge3_12_3"%string, 9)) [(EVar "_60"%string);(EVar "_61"%string);(EVar "_62"%string);(EVar "_63"%string);(EVar "_64"%string);(EVar "_65"%string);(EVar "_66"%string);(ECons (EVar "_67"%string) (EVar "_69"%string));(EVar "_68"%string)]))]));([(PVar "E1"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "E2"%string);(EVar "HdM"%string)]), (EApp (EFunId ("ukeymerge3_2"%string, 11)) [(EVar "I"%string);(EVar "E1"%string);(EVar "T1"%string);(EVar "H1"%string);(EVar "T2"%string);(EVar "HdM"%string);(EVar "T2"%string);(EVar "M"%string);(EVar "E3"%string);(EVar "H3"%string);(EVar "T3"%string)]));([(PVar "E1"%string)], (ELit (Atom "true"%string)), (ECase (EValues [(EVar "I"%string);(EVar "E1"%string);(EVar "T1"%string);(EVar "H1"%string);(EVar "E2"%string);(EVar "H2"%string);(EVar "T2"%string);(EVar "E3"%string);(EVar "H3"%string);(EVar "T3"%string);(EVar "M"%string);(EVar "HdM"%string);(EVar "T2"%string)]) [([(PVar "_81"%string);(PVar "_82"%string);(PVar "_83"%string);(PVar "_84"%string);(PVar "_85"%string);(PVar "_86"%string);(PVar "_87"%string);(PVar "_88"%string);(PVar "_89"%string);(PVar "_90"%string);(PVar "_91"%string);(PVar "_HdM"%string);(PVar "_92"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "_85"%string);(EVar "_88"%string)]), (EApp (EFunId ("ukeymerge3_2"%string, 11)) [(EVar "_81"%string);(EVar "_82"%string);(EVar "_83"%string);(EVar "_84"%string);(EVar "_87"%string);(EVar "_85"%string);(EVar "_92"%string);(ECons (EVar "_86"%string) (EVar "_91"%string));(EVar "_88"%string);(EVar "_89"%string);(EVar "_90"%string)]));([(PVar "_93"%string);(PVar "_94"%string);(PVar "_95"%string);(PVar "_96"%string);(PVar "_97"%string);(PVar "_98"%string);(PVar "_99"%string);(PVar "_100"%string);(PVar "_H3"%string);(PVar "_101"%string);(PVar "_102"%string);(PVar "_103"%string);(PVar "_D"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "_100"%string);(EVar "_103"%string)]), (EApp (EFunId ("ukeymerge3_21_3"%string, 9)) [(EVar "_93"%string);(EVar "_94"%string);(EVar "_95"%string);(EVar "_96"%string);(EVar "_97"%string);(EVar "_98"%string);(EVar "_99"%string);(EVar "_102"%string);(EVar "_101"%string)]));([(PVar "_104"%string);(PVar "_105"%string);(PVar "_106"%string);(PVar "_107"%string);(PVar "_108"%string);(PVar "_109"%string);(PVar "_110"%string);(PVar "_E3"%string);(PVar "_111"%string);(PVar "_112"%string);(PVar "_113"%string);(PVar "_HdM"%string);(PVar "_D"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("ukeymerge3_21_3"%string, 9)) [(EVar "_104"%string);(EVar "_105"%string);(EVar "_106"%string);(EVar "_107"%string);(EVar "_108"%string);(EVar "_109"%string);(EVar "_110"%string);(ECons (EVar "_111"%string) (EVar "_113"%string));(EVar "_112"%string)]))]))]));([(PVar "I"%string);PNil;(PVar "_D"%string);(PVar "HdM"%string);(PVar "E2"%string);(PVar "_H2"%string);(PVar "T2"%string);(PVar "M"%string);(PVar "E3"%string);(PVar "H3"%string);(PVar "T3"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "E2"%string);(EVar "HdM"%string)]), (EApp (EFunId ("ukeymerge2_1"%string, 7)) [(EVar "I"%string);(EVar "T2"%string);(EVar "E3"%string);(EVar "HdM"%string);(EVar "T3"%string);(EVar "M"%string);(EVar "H3"%string)]));([(PVar "I"%string);PNil;(PVar "_D"%string);(PVar "_HdM"%string);(PVar "E2"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "M"%string);(PVar "E3"%string);(PVar "H3"%string);(PVar "T3"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "E2"%string);(EVar "E3"%string)]), (EApp (EFunId ("ukeymerge2_1"%string, 7)) [(EVar "I"%string);(EVar "T2"%string);(EVar "E3"%string);(EVar "E2"%string);(EVar "T3"%string);(ECons (EVar "H2"%string) (EVar "M"%string));(EVar "H3"%string)]));([(PVar "I"%string);PNil;(PVar "_D"%string);(PVar "HdM"%string);(PVar "E2"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "M"%string);(PVar "E3"%string);(PVar "_H3"%string);(PVar "T3"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "E3"%string);(EVar "HdM"%string)]), (EApp (EFunId ("ukeymerge2_2"%string, 6)) [(EVar "I"%string);(EVar "T2"%string);(EVar "E2"%string);(EVar "H2"%string);(EVar "T3"%string);(EVar "M"%string)]));([(PVar "I"%string);PNil;(PVar "_D"%string);(PVar "_HdM"%string);(PVar "E2"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "M"%string);(PVar "_E3"%string);(PVar "H3"%string);(PVar "T3"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("ukeymerge2_2"%string, 6)) [(EVar "I"%string);(EVar "T2"%string);(EVar "E2"%string);(EVar "H2"%string);(EVar "T3"%string);(ECons (EVar "H3"%string) (EVar "M"%string))]));([(PVar "_22"%string);(PVar "_21"%string);(PVar "_20"%string);(PVar "_19"%string);(PVar "_18"%string);(PVar "_17"%string);(PVar "_16"%string);(PVar "_15"%string);(PVar "_14"%string);(PVar "_13"%string);(PVar "_12"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_22"%string);(EVar "_21"%string);(EVar "_20"%string);(EVar "_19"%string);(EVar "_18"%string);(EVar "_17"%string);(EVar "_16"%string);(EVar "_15"%string);(EVar "_14"%string);(EVar "_13"%string);(EVar "_12"%string)])]))]) |};
          {| identifier := ("ukeymerge3_2"%string, 11) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string;"_6"%string;"_7"%string;"_8"%string;"_9"%string;"_10"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string);(EVar "_6"%string);(EVar "_7"%string);(EVar "_8"%string);(EVar "_9"%string);(EVar "_10"%string)]) [([(PVar "I"%string);(PVar "E1"%string);(PVar "T1"%string);(PVar "H1"%string);(PCons (PVar "H2"%string) (PVar "T2"%string));(PVar "HdM"%string);(PVar "D"%string);(PVar "M"%string);(PVar "E3"%string);(PVar "H3"%string);(PVar "T3"%string)], (ELit (Atom "true"%string)), (ECase (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "I"%string);(EVar "H2"%string)]) [([(PVar "E2"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "E1"%string);(EVar "E2"%string)]), (ECase (EValues [(EVar "I"%string);(EVar "E1"%string);(EVar "T1"%string);(EVar "H1"%string);(EVar "E2"%string);(EVar "H2"%string);(EVar "T2"%string);(EVar "E3"%string);(EVar "H3"%string);(EVar "T3"%string);(EVar "M"%string);(EVar "HdM"%string);(EVar "T1"%string)]) [([(PVar "_37"%string);(PVar "_38"%string);(PVar "_39"%string);(PVar "_40"%string);(PVar "_41"%string);(PVar "_42"%string);(PVar "_43"%string);(PVar "_44"%string);(PVar "_45"%string);(PVar "_46"%string);(PVar "_47"%string);(PVar "_HdM"%string);(PVar "_48"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "_38"%string);(EVar "_44"%string)]), (EApp (EFunId ("ukeymerge3_1"%string, 11)) [(EVar "_37"%string);(EVar "_39"%string);(EVar "_48"%string);(EVar "_38"%string);(EVar "_41"%string);(EVar "_42"%string);(EVar "_43"%string);(ECons (EVar "_40"%string) (EVar "_47"%string));(EVar "_44"%string);(EVar "_45"%string);(EVar "_46"%string)]));([(PVar "_49"%string);(PVar "_50"%string);(PVar "_51"%string);(PVar "_52"%string);(PVar "_53"%string);(PVar "_54"%string);(PVar "_55"%string);(PVar "_56"%string);(PVar "_H3"%string);(PVar "_57"%string);(PVar "_58"%string);(PVar "_59"%string);(PVar "_D"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "_56"%string);(EVar "_59"%string)]), (EApp (EFunId ("ukeymerge3_12_3"%string, 9)) [(EVar "_49"%string);(EVar "_50"%string);(EVar "_51"%string);(EVar "_52"%string);(EVar "_53"%string);(EVar "_54"%string);(EVar "_55"%string);(EVar "_58"%string);(EVar "_57"%string)]));([(PVar "_60"%string);(PVar "_61"%string);(PVar "_62"%string);(PVar "_63"%string);(PVar "_64"%string);(PVar "_65"%string);(PVar "_66"%string);(PVar "_E3"%string);(PVar "_67"%string);(PVar "_68"%string);(PVar "_69"%string);(PVar "_HdM"%string);(PVar "_D"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("ukeymerge3_12_3"%string, 9)) [(EVar "_60"%string);(EVar "_61"%string);(EVar "_62"%string);(EVar "_63"%string);(EVar "_64"%string);(EVar "_65"%string);(EVar "_66"%string);(ECons (EVar "_67"%string) (EVar "_69"%string));(EVar "_68"%string)]))]));([(PVar "E2"%string)], (ELit (Atom "true"%string)), (ECase (EValues [(EVar "I"%string);(EVar "E1"%string);(EVar "T1"%string);(EVar "H1"%string);(EVar "E2"%string);(EVar "H2"%string);(EVar "T2"%string);(EVar "E3"%string);(EVar "H3"%string);(EVar "T3"%string);(EVar "M"%string);(EVar "HdM"%string);(EVar "D"%string)]) [([(PVar "_81"%string);(PVar "_82"%string);(PVar "_83"%string);(PVar "_84"%string);(PVar "_85"%string);(PVar "_86"%string);(PVar "_87"%string);(PVar "_88"%string);(PVar "_89"%string);(PVar "_90"%string);(PVar "_91"%string);(PVar "_HdM"%string);(PVar "_92"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "_85"%string);(EVar "_88"%string)]), (EApp (EFunId ("ukeymerge3_2"%string, 11)) [(EVar "_81"%string);(EVar "_82"%string);(EVar "_83"%string);(EVar "_84"%string);(EVar "_87"%string);(EVar "_85"%string);(EVar "_92"%string);(ECons (EVar "_86"%string) (EVar "_91"%string));(EVar "_88"%string);(EVar "_89"%string);(EVar "_90"%string)]));([(PVar "_93"%string);(PVar "_94"%string);(PVar "_95"%string);(PVar "_96"%string);(PVar "_97"%string);(PVar "_98"%string);(PVar "_99"%string);(PVar "_100"%string);(PVar "_H3"%string);(PVar "_101"%string);(PVar "_102"%string);(PVar "_103"%string);(PVar "_D"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "_100"%string);(EVar "_103"%string)]), (EApp (EFunId ("ukeymerge3_21_3"%string, 9)) [(EVar "_93"%string);(EVar "_94"%string);(EVar "_95"%string);(EVar "_96"%string);(EVar "_97"%string);(EVar "_98"%string);(EVar "_99"%string);(EVar "_102"%string);(EVar "_101"%string)]));([(PVar "_104"%string);(PVar "_105"%string);(PVar "_106"%string);(PVar "_107"%string);(PVar "_108"%string);(PVar "_109"%string);(PVar "_110"%string);(PVar "_E3"%string);(PVar "_111"%string);(PVar "_112"%string);(PVar "_113"%string);(PVar "_HdM"%string);(PVar "_D"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("ukeymerge3_21_3"%string, 9)) [(EVar "_104"%string);(EVar "_105"%string);(EVar "_106"%string);(EVar "_107"%string);(EVar "_108"%string);(EVar "_109"%string);(EVar "_110"%string);(ECons (EVar "_111"%string) (EVar "_113"%string));(EVar "_112"%string)]))]))]));([(PVar "I"%string);(PVar "E1"%string);(PVar "T1"%string);(PVar "H1"%string);PNil;(PVar "_HdM"%string);(PVar "_D"%string);(PVar "M"%string);(PVar "E3"%string);(PVar "H3"%string);(PVar "T3"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "E1"%string);(EVar "E3"%string)]), (EApp (EFunId ("ukeymerge2_1"%string, 7)) [(EVar "I"%string);(EVar "T1"%string);(EVar "E3"%string);(EVar "E1"%string);(EVar "T3"%string);(ECons (EVar "H1"%string) (EVar "M"%string));(EVar "H3"%string)]));([(PVar "I"%string);(PVar "E1"%string);(PVar "T1"%string);(PVar "H1"%string);PNil;(PVar "HdM"%string);(PVar "_D"%string);(PVar "M"%string);(PVar "E3"%string);(PVar "_H3"%string);(PVar "T3"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "E3"%string);(EVar "HdM"%string)]), (EApp (EFunId ("ukeymerge2_2"%string, 6)) [(EVar "I"%string);(EVar "T1"%string);(EVar "E1"%string);(EVar "H1"%string);(EVar "T3"%string);(EVar "M"%string)]));([(PVar "I"%string);(PVar "E1"%string);(PVar "T1"%string);(PVar "H1"%string);PNil;(PVar "_HdM"%string);(PVar "_D"%string);(PVar "M"%string);(PVar "_E3"%string);(PVar "H3"%string);(PVar "T3"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("ukeymerge2_2"%string, 6)) [(EVar "I"%string);(EVar "T1"%string);(EVar "E1"%string);(EVar "H1"%string);(EVar "T3"%string);(ECons (EVar "H3"%string) (EVar "M"%string))]));([(PVar "_22"%string);(PVar "_21"%string);(PVar "_20"%string);(PVar "_19"%string);(PVar "_18"%string);(PVar "_17"%string);(PVar "_16"%string);(PVar "_15"%string);(PVar "_14"%string);(PVar "_13"%string);(PVar "_12"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_22"%string);(EVar "_21"%string);(EVar "_20"%string);(EVar "_19"%string);(EVar "_18"%string);(EVar "_17"%string);(EVar "_16"%string);(EVar "_15"%string);(EVar "_14"%string);(EVar "_13"%string);(EVar "_12"%string)])]))]) |};
          {| identifier := ("ukeymerge3_12"%string, 13) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string;"_6"%string;"_7"%string;"_8"%string;"_9"%string;"_10"%string;"_11"%string;"_12"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string);(EVar "_6"%string);(EVar "_7"%string);(EVar "_8"%string);(EVar "_9"%string);(EVar "_10"%string);(EVar "_11"%string);(EVar "_12"%string)]) [([(PVar "I"%string);(PVar "E1"%string);(PVar "T1"%string);(PVar "H1"%string);(PVar "E2"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "E3"%string);(PVar "H3"%string);(PVar "T3"%string);(PVar "M"%string);(PVar "_HdM"%string);(PVar "D"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "E1"%string);(EVar "E3"%string)]), (EApp (EFunId ("ukeymerge3_1"%string, 11)) [(EVar "I"%string);(EVar "T1"%string);(EVar "D"%string);(EVar "E1"%string);(EVar "E2"%string);(EVar "H2"%string);(EVar "T2"%string);(ECons (EVar "H1"%string) (EVar "M"%string));(EVar "E3"%string);(EVar "H3"%string);(EVar "T3"%string)]));([(PVar "I"%string);(PVar "E1"%string);(PVar "T1"%string);(PVar "H1"%string);(PVar "E2"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "E3"%string);(PVar "_H3"%string);(PVar "T3"%string);(PVar "M"%string);(PVar "HdM"%string);(PVar "_D"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "E3"%string);(EVar "HdM"%string)]), (EApp (EFunId ("ukeymerge3_12_3"%string, 9)) [(EVar "I"%string);(EVar "E1"%string);(EVar "T1"%string);(EVar "H1"%string);(EVar "E2"%string);(EVar "H2"%string);(EVar "T2"%string);(EVar "M"%string);(EVar "T3"%string)]));([(PVar "I"%string);(PVar "E1"%string);(PVar "T1"%string);(PVar "H1"%string);(PVar "E2"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "_E3"%string);(PVar "H3"%string);(PVar "T3"%string);(PVar "M"%string);(PVar "_HdM"%string);(PVar "_D"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("ukeymerge3_12_3"%string, 9)) [(EVar "I"%string);(EVar "E1"%string);(EVar "T1"%string);(EVar "H1"%string);(EVar "E2"%string);(EVar "H2"%string);(EVar "T2"%string);(ECons (EVar "H3"%string) (EVar "M"%string));(EVar "T3"%string)]))]) |};
          {| identifier := ("ukeymerge3_12_3"%string, 9) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string;"_6"%string;"_7"%string;"_8"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string);(EVar "_6"%string);(EVar "_7"%string);(EVar "_8"%string)]) [([(PVar "I"%string);(PVar "E1"%string);(PVar "T1"%string);(PVar "H1"%string);(PVar "E2"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "M"%string);(PCons (PVar "H3"%string) (PVar "T3"%string))], (ELit (Atom "true"%string)), (ECase (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "I"%string);(EVar "H3"%string)]) [([(PVar "E3"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "E1"%string);(EVar "E3"%string)]), (EApp (EFunId ("ukeymerge3_1"%string, 11)) [(EVar "I"%string);(EVar "T1"%string);(EVar "T1"%string);(EVar "E1"%string);(EVar "E2"%string);(EVar "H2"%string);(EVar "T2"%string);(ECons (EVar "H1"%string) (EVar "M"%string));(EVar "E3"%string);(EVar "H3"%string);(EVar "T3"%string)]));([(PVar "_E3"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("ukeymerge3_12_3"%string, 9)) [(EVar "I"%string);(EVar "E1"%string);(EVar "T1"%string);(EVar "H1"%string);(EVar "E2"%string);(EVar "H2"%string);(EVar "T2"%string);(ECons (EVar "H3"%string) (EVar "M"%string));(EVar "T3"%string)]))]));([(PVar "I"%string);(PVar "E1"%string);(PVar "T1"%string);(PVar "H1"%string);(PVar "E2"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "M"%string);PNil], (ELit (Atom "true"%string)), (EApp (EFunId ("ukeymerge2_1"%string, 7)) [(EVar "I"%string);(EVar "T1"%string);(EVar "E2"%string);(EVar "E1"%string);(EVar "T2"%string);(ECons (EVar "H1"%string) (EVar "M"%string));(EVar "H2"%string)]));([(PVar "_18"%string);(PVar "_17"%string);(PVar "_16"%string);(PVar "_15"%string);(PVar "_14"%string);(PVar "_13"%string);(PVar "_12"%string);(PVar "_11"%string);(PVar "_10"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_18"%string);(EVar "_17"%string);(EVar "_16"%string);(EVar "_15"%string);(EVar "_14"%string);(EVar "_13"%string);(EVar "_12"%string);(EVar "_11"%string);(EVar "_10"%string)])]))]) |};
          {| identifier := ("ukeymerge3_21"%string, 13) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string;"_6"%string;"_7"%string;"_8"%string;"_9"%string;"_10"%string;"_11"%string;"_12"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string);(EVar "_6"%string);(EVar "_7"%string);(EVar "_8"%string);(EVar "_9"%string);(EVar "_10"%string);(EVar "_11"%string);(EVar "_12"%string)]) [([(PVar "I"%string);(PVar "E1"%string);(PVar "T1"%string);(PVar "H1"%string);(PVar "E2"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "E3"%string);(PVar "H3"%string);(PVar "T3"%string);(PVar "M"%string);(PVar "_HdM"%string);(PVar "D"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "E2"%string);(EVar "E3"%string)]), (EApp (EFunId ("ukeymerge3_2"%string, 11)) [(EVar "I"%string);(EVar "E1"%string);(EVar "T1"%string);(EVar "H1"%string);(EVar "T2"%string);(EVar "E2"%string);(EVar "D"%string);(ECons (EVar "H2"%string) (EVar "M"%string));(EVar "E3"%string);(EVar "H3"%string);(EVar "T3"%string)]));([(PVar "I"%string);(PVar "E1"%string);(PVar "T1"%string);(PVar "H1"%string);(PVar "E2"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "E3"%string);(PVar "_H3"%string);(PVar "T3"%string);(PVar "M"%string);(PVar "HdM"%string);(PVar "_D"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "E3"%string);(EVar "HdM"%string)]), (EApp (EFunId ("ukeymerge3_21_3"%string, 9)) [(EVar "I"%string);(EVar "E1"%string);(EVar "T1"%string);(EVar "H1"%string);(EVar "E2"%string);(EVar "H2"%string);(EVar "T2"%string);(EVar "M"%string);(EVar "T3"%string)]));([(PVar "I"%string);(PVar "E1"%string);(PVar "T1"%string);(PVar "H1"%string);(PVar "E2"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "_E3"%string);(PVar "H3"%string);(PVar "T3"%string);(PVar "M"%string);(PVar "_HdM"%string);(PVar "_D"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("ukeymerge3_21_3"%string, 9)) [(EVar "I"%string);(EVar "E1"%string);(EVar "T1"%string);(EVar "H1"%string);(EVar "E2"%string);(EVar "H2"%string);(EVar "T2"%string);(ECons (EVar "H3"%string) (EVar "M"%string));(EVar "T3"%string)]))]) |};
          {| identifier := ("ukeymerge3_21_3"%string, 9) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string;"_6"%string;"_7"%string;"_8"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string);(EVar "_6"%string);(EVar "_7"%string);(EVar "_8"%string)]) [([(PVar "I"%string);(PVar "E1"%string);(PVar "T1"%string);(PVar "H1"%string);(PVar "E2"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "M"%string);(PCons (PVar "H3"%string) (PVar "T3"%string))], (ELit (Atom "true"%string)), (ECase (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "I"%string);(EVar "H3"%string)]) [([(PVar "E3"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "E2"%string);(EVar "E3"%string)]), (EApp (EFunId ("ukeymerge3_2"%string, 11)) [(EVar "I"%string);(EVar "E1"%string);(EVar "T1"%string);(EVar "H1"%string);(EVar "T2"%string);(EVar "E2"%string);(EVar "T2"%string);(ECons (EVar "H2"%string) (EVar "M"%string));(EVar "E3"%string);(EVar "H3"%string);(EVar "T3"%string)]));([(PVar "_E3"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("ukeymerge3_21_3"%string, 9)) [(EVar "I"%string);(EVar "E1"%string);(EVar "T1"%string);(EVar "H1"%string);(EVar "E2"%string);(EVar "H2"%string);(EVar "T2"%string);(ECons (EVar "H3"%string) (EVar "M"%string));(EVar "T3"%string)]))]));([(PVar "I"%string);(PVar "E1"%string);(PVar "T1"%string);(PVar "H1"%string);(PVar "_E2"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "M"%string);PNil], (ELit (Atom "true"%string)), (EApp (EFunId ("ukeymerge2_2"%string, 6)) [(EVar "I"%string);(EVar "T1"%string);(EVar "E1"%string);(EVar "H1"%string);(EVar "T2"%string);(ECons (EVar "H2"%string) (EVar "M"%string))]));([(PVar "_18"%string);(PVar "_17"%string);(PVar "_16"%string);(PVar "_15"%string);(PVar "_14"%string);(PVar "_13"%string);(PVar "_12"%string);(PVar "_11"%string);(PVar "_10"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_18"%string);(EVar "_17"%string);(EVar "_16"%string);(EVar "_15"%string);(EVar "_14"%string);(EVar "_13"%string);(EVar "_12"%string);(EVar "_11"%string);(EVar "_10"%string)])]))]) |};
          {| identifier := ("rukeymerge3_1"%string, 11) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string;"_6"%string;"_7"%string;"_8"%string;"_9"%string;"_10"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string);(EVar "_6"%string);(EVar "_7"%string);(EVar "_8"%string);(EVar "_9"%string);(EVar "_10"%string)]) [([(PVar "I"%string);(PCons (PVar "H1"%string) (PVar "T1"%string));(PVar "D1"%string);(PVar "D2"%string);(PVar "E2"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "M"%string);(PVar "E3"%string);(PVar "H3"%string);(PVar "T3"%string)], (ELit (Atom "true"%string)), (ECase (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "I"%string);(EVar "H1"%string)]) [([(PVar "E1"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "E1"%string);(EVar "E2"%string)]), (ECase (EValues [(EVar "I"%string);(EVar "E1"%string);(EVar "H1"%string);(EVar "T1"%string);(EVar "E2"%string);(EVar "H2"%string);(EVar "T2"%string);(EVar "E3"%string);(EVar "H3"%string);(EVar "T3"%string);(EVar "M"%string)]) [([(PVar "_37"%string);(PVar "_38"%string);(PVar "_39"%string);(PVar "_40"%string);(PVar "_41"%string);(PVar "_42"%string);(PVar "_43"%string);(PVar "_44"%string);(PVar "_45"%string);(PVar "_46"%string);(PVar "_47"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "_41"%string);(EVar "_44"%string)]), (EApp (EFunId ("rukeymerge3_12_3"%string, 11)) [(EVar "_37"%string);(EVar "_38"%string);(EVar "_39"%string);(EVar "_40"%string);(EVar "_41"%string);(EVar "_42"%string);(EVar "_43"%string);(EVar "_47"%string);(EVar "_44"%string);(EVar "_45"%string);(EVar "_46"%string)]));([(PVar "_48"%string);(PVar "_49"%string);(PVar "_50"%string);(PVar "_51"%string);(PVar "_52"%string);(PVar "_53"%string);(PVar "_54"%string);(PVar "_55"%string);(PVar "_56"%string);(PVar "_57"%string);(PVar "_58"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rukeymerge3_2"%string, 11)) [(EVar "_48"%string);(EVar "_49"%string);(EVar "_50"%string);(EVar "_51"%string);(EVar "_54"%string);(EVar "_53"%string);(EVar "_52"%string);(EVar "_58"%string);(EVar "_55"%string);(EVar "_56"%string);(EVar "_57"%string)]))]));([(PVar "E1"%string)], (ELit (Atom "true"%string)), (ECase (EValues [(EVar "I"%string);(EVar "E1"%string);(EVar "H1"%string);(EVar "T1"%string);(EVar "E2"%string);(EVar "H2"%string);(EVar "T2"%string);(EVar "E3"%string);(EVar "H3"%string);(EVar "T3"%string);(EVar "M"%string);(EVar "D1"%string);(EVar "D2"%string)]) [([(PVar "_70"%string);(PVar "_71"%string);(PVar "_72"%string);(PVar "_73"%string);(PVar "_74"%string);(PVar "_75"%string);(PVar "_76"%string);(PVar "_77"%string);(PVar "_78"%string);(PVar "_79"%string);(PVar "_80"%string);(PVar "_D1"%string);(PVar "_D2"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "_71"%string);(EVar "_77"%string)]), (EApp (EFunId ("rukeymerge3_21_3"%string, 11)) [(EVar "_70"%string);(EVar "_71"%string);(EVar "_72"%string);(EVar "_73"%string);(EVar "_74"%string);(EVar "_75"%string);(EVar "_76"%string);(EVar "_80"%string);(EVar "_77"%string);(EVar "_78"%string);(EVar "_79"%string)]));([(PVar "_81"%string);(PVar "_E1"%string);(PVar "_82"%string);(PVar "_83"%string);(PVar "_84"%string);(PVar "_85"%string);(PVar "_86"%string);(PVar "_87"%string);(PVar "_88"%string);(PVar "_89"%string);(PVar "_90"%string);(PVar "_91"%string);(PVar "_92"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rukeymerge3_1"%string, 11)) [(EVar "_81"%string);(EVar "_83"%string);(EVar "_91"%string);(EVar "_92"%string);(EVar "_84"%string);(EVar "_85"%string);(EVar "_86"%string);(ECons (EVar "_82"%string) (EVar "_90"%string));(EVar "_87"%string);(EVar "_88"%string);(EVar "_89"%string)]))]))]));([(PVar "I"%string);PNil;(PVar "_D1"%string);(PVar "_D2"%string);(PVar "E2"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "M"%string);(PVar "E3"%string);(PVar "H3"%string);(PVar "T3"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "E2"%string);(EVar "E3"%string)]), (EApp (EFunId ("rukeymerge2_2"%string, 8)) [(EVar "I"%string);(EVar "T2"%string);(EVar "E2"%string);(EVar "T3"%string);(EVar "M"%string);(EVar "E3"%string);(EVar "H3"%string);(EVar "H2"%string)]));([(PVar "I"%string);PNil;(PVar "_D1"%string);(PVar "_D2"%string);(PVar "_E2"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "M"%string);(PVar "E3"%string);(PVar "H3"%string);(PVar "T3"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rukeymerge2_1"%string, 6)) [(EVar "I"%string);(EVar "T2"%string);(EVar "E3"%string);(EVar "T3"%string);(ECons (EVar "H2"%string) (EVar "M"%string));(EVar "H3"%string)]));([(PVar "_22"%string);(PVar "_21"%string);(PVar "_20"%string);(PVar "_19"%string);(PVar "_18"%string);(PVar "_17"%string);(PVar "_16"%string);(PVar "_15"%string);(PVar "_14"%string);(PVar "_13"%string);(PVar "_12"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_22"%string);(EVar "_21"%string);(EVar "_20"%string);(EVar "_19"%string);(EVar "_18"%string);(EVar "_17"%string);(EVar "_16"%string);(EVar "_15"%string);(EVar "_14"%string);(EVar "_13"%string);(EVar "_12"%string)])]))]) |};
          {| identifier := ("rukeymerge3_12a"%string, 11) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string;"_6"%string;"_7"%string;"_8"%string;"_9"%string;"_10"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string);(EVar "_6"%string);(EVar "_7"%string);(EVar "_8"%string);(EVar "_9"%string);(EVar "_10"%string)]) [([(PVar "I"%string);(PVar "E1"%string);(PVar "H1"%string);(PVar "T1"%string);(PVar "E2"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "E3"%string);(PVar "H3"%string);(PVar "T3"%string);(PVar "M"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "E2"%string);(EVar "E3"%string)]), (EApp (EFunId ("rukeymerge3_12_3"%string, 11)) [(EVar "I"%string);(EVar "E1"%string);(EVar "H1"%string);(EVar "T1"%string);(EVar "E2"%string);(EVar "H2"%string);(EVar "T2"%string);(EVar "M"%string);(EVar "E3"%string);(EVar "H3"%string);(EVar "T3"%string)]));([(PVar "I"%string);(PVar "E1"%string);(PVar "H1"%string);(PVar "T1"%string);(PVar "E2"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "E3"%string);(PVar "H3"%string);(PVar "T3"%string);(PVar "M"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rukeymerge3_2"%string, 11)) [(EVar "I"%string);(EVar "E1"%string);(EVar "H1"%string);(EVar "T1"%string);(EVar "T2"%string);(EVar "H2"%string);(EVar "E2"%string);(EVar "M"%string);(EVar "E3"%string);(EVar "H3"%string);(EVar "T3"%string)]))]) |};
          {| identifier := ("rukeymerge3_21a"%string, 13) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string;"_6"%string;"_7"%string;"_8"%string;"_9"%string;"_10"%string;"_11"%string;"_12"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string);(EVar "_6"%string);(EVar "_7"%string);(EVar "_8"%string);(EVar "_9"%string);(EVar "_10"%string);(EVar "_11"%string);(EVar "_12"%string)]) [([(PVar "I"%string);(PVar "E1"%string);(PVar "H1"%string);(PVar "T1"%string);(PVar "E2"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "E3"%string);(PVar "H3"%string);(PVar "T3"%string);(PVar "M"%string);(PVar "_D1"%string);(PVar "_D2"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "E1"%string);(EVar "E3"%string)]), (EApp (EFunId ("rukeymerge3_21_3"%string, 11)) [(EVar "I"%string);(EVar "E1"%string);(EVar "H1"%string);(EVar "T1"%string);(EVar "E2"%string);(EVar "H2"%string);(EVar "T2"%string);(EVar "M"%string);(EVar "E3"%string);(EVar "H3"%string);(EVar "T3"%string)]));([(PVar "I"%string);(PVar "_E1"%string);(PVar "H1"%string);(PVar "T1"%string);(PVar "E2"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "E3"%string);(PVar "H3"%string);(PVar "T3"%string);(PVar "M"%string);(PVar "D1"%string);(PVar "D2"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rukeymerge3_1"%string, 11)) [(EVar "I"%string);(EVar "T1"%string);(EVar "D1"%string);(EVar "D2"%string);(EVar "E2"%string);(EVar "H2"%string);(EVar "T2"%string);(ECons (EVar "H1"%string) (EVar "M"%string));(EVar "E3"%string);(EVar "H3"%string);(EVar "T3"%string)]))]) |};
          {| identifier := ("rukeymerge3_2"%string, 11) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string;"_6"%string;"_7"%string;"_8"%string;"_9"%string;"_10"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string);(EVar "_6"%string);(EVar "_7"%string);(EVar "_8"%string);(EVar "_9"%string);(EVar "_10"%string)]) [([(PVar "I"%string);(PVar "E1"%string);(PVar "H1"%string);(PVar "T1"%string);(PCons (PVar "H2"%string) (PVar "T2"%string));(PVar "H2M"%string);(PVar "E2M"%string);(PVar "M"%string);(PVar "E3"%string);(PVar "H3"%string);(PVar "T3"%string)], (ELit (Atom "true"%string)), (ECase (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "I"%string);(EVar "H2"%string)]) [([(PVar "E2"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "E1"%string);(EVar "E2"%string)]), (ECase (EValues [(EVar "I"%string);(EVar "E1"%string);(EVar "H1"%string);(EVar "T1"%string);(EVar "E2"%string);(EVar "H2"%string);(EVar "T2"%string);(EVar "E3"%string);(EVar "H3"%string);(EVar "T3"%string);(EVar "M"%string);(EVar "H2M"%string)]) [([(PVar "_35"%string);(PVar "_36"%string);(PVar "_37"%string);(PVar "_38"%string);(PVar "_39"%string);(PVar "_40"%string);(PVar "_41"%string);(PVar "_42"%string);(PVar "_43"%string);(PVar "_44"%string);(PVar "_45"%string);(PVar "_46"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "_39"%string);(EVar "_42"%string)]), (EApp (EFunId ("rukeymerge3_12_3"%string, 11)) [(EVar "_35"%string);(EVar "_36"%string);(EVar "_37"%string);(EVar "_38"%string);(EVar "_39"%string);(EVar "_40"%string);(EVar "_41"%string);(ECons (EVar "_46"%string) (EVar "_45"%string));(EVar "_42"%string);(EVar "_43"%string);(EVar "_44"%string)]));([(PVar "_47"%string);(PVar "_48"%string);(PVar "_49"%string);(PVar "_50"%string);(PVar "_51"%string);(PVar "_52"%string);(PVar "_53"%string);(PVar "_54"%string);(PVar "_55"%string);(PVar "_56"%string);(PVar "_57"%string);(PVar "_58"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rukeymerge3_2"%string, 11)) [(EVar "_47"%string);(EVar "_48"%string);(EVar "_49"%string);(EVar "_50"%string);(EVar "_53"%string);(EVar "_52"%string);(EVar "_51"%string);(ECons (EVar "_58"%string) (EVar "_57"%string));(EVar "_54"%string);(EVar "_55"%string);(EVar "_56"%string)]))]));([(PVar "E2"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "E1"%string);(EVar "E2M"%string)]), (EApp (EFunId ("rukeymerge3_1"%string, 11)) [(EVar "I"%string);(EVar "T1"%string);(EVar "H1"%string);(EVar "T1"%string);(EVar "E2"%string);(EVar "H2"%string);(EVar "T2"%string);(ECons (EVar "H1"%string) (EVar "M"%string));(EVar "E3"%string);(EVar "H3"%string);(EVar "T3"%string)]));([(PVar "E2"%string)], (ELit (Atom "true"%string)), (ECase (EValues [(EVar "I"%string);(EVar "E1"%string);(EVar "H1"%string);(EVar "T1"%string);(EVar "E2"%string);(EVar "H2"%string);(EVar "T2"%string);(EVar "E3"%string);(EVar "H3"%string);(EVar "T3"%string);(EVar "M"%string);(EVar "H2M"%string)]) [([(PVar "_70"%string);(PVar "_71"%string);(PVar "_72"%string);(PVar "_73"%string);(PVar "_74"%string);(PVar "_75"%string);(PVar "_76"%string);(PVar "_77"%string);(PVar "_78"%string);(PVar "_79"%string);(PVar "_80"%string);(PVar "_81"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "_71"%string);(EVar "_77"%string)]), (EApp (EFunId ("rukeymerge3_21_3"%string, 11)) [(EVar "_70"%string);(EVar "_71"%string);(EVar "_72"%string);(EVar "_73"%string);(EVar "_74"%string);(EVar "_75"%string);(EVar "_76"%string);(ECons (EVar "_81"%string) (EVar "_80"%string));(EVar "_77"%string);(EVar "_78"%string);(EVar "_79"%string)]));([(PVar "_82"%string);(PVar "_E1"%string);(PVar "_83"%string);(PVar "_84"%string);(PVar "_85"%string);(PVar "_86"%string);(PVar "_87"%string);(PVar "_88"%string);(PVar "_89"%string);(PVar "_90"%string);(PVar "_91"%string);(PVar "_92"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rukeymerge3_1"%string, 11)) [(EVar "_82"%string);(EVar "_84"%string);(EVar "_83"%string);(EVar "_84"%string);(EVar "_85"%string);(EVar "_86"%string);(EVar "_87"%string);(ECons (EVar "_83"%string) (ECons (EVar "_92"%string) (EVar "_91"%string)));(EVar "_88"%string);(EVar "_89"%string);(EVar "_90"%string)]))]))]));([(PVar "I"%string);(PVar "E1"%string);(PVar "H1"%string);(PVar "T1"%string);PNil;(PVar "_H2M"%string);(PVar "E2M"%string);(PVar "M"%string);(PVar "E3"%string);(PVar "H3"%string);(PVar "T3"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "E1"%string);(EVar "E2M"%string)]), (EApp (EFunId ("rukeymerge2_1"%string, 6)) [(EVar "I"%string);(EVar "T1"%string);(EVar "E3"%string);(EVar "T3"%string);(ECons (EVar "H1"%string) (EVar "M"%string));(EVar "H3"%string)]));([(PVar "I"%string);(PVar "E1"%string);(PVar "H1"%string);(PVar "T1"%string);PNil;(PVar "H2M"%string);(PVar "_E2M"%string);(PVar "M"%string);(PVar "E3"%string);(PVar "H3"%string);(PVar "T3"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "E1"%string);(EVar "E3"%string)]), (EApp (EFunId ("rukeymerge2_2"%string, 8)) [(EVar "I"%string);(EVar "T1"%string);(EVar "E1"%string);(EVar "T3"%string);(ECons (EVar "H2M"%string) (EVar "M"%string));(EVar "E3"%string);(EVar "H3"%string);(EVar "H1"%string)]));([(PVar "I"%string);(PVar "_E1"%string);(PVar "H1"%string);(PVar "T1"%string);PNil;(PVar "H2M"%string);(PVar "_E2M"%string);(PVar "M"%string);(PVar "E3"%string);(PVar "H3"%string);(PVar "T3"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rukeymerge2_1"%string, 6)) [(EVar "I"%string);(EVar "T1"%string);(EVar "E3"%string);(EVar "T3"%string);(ECons (EVar "H1"%string) (ECons (EVar "H2M"%string) (EVar "M"%string)));(EVar "H3"%string)]));([(PVar "_22"%string);(PVar "_21"%string);(PVar "_20"%string);(PVar "_19"%string);(PVar "_18"%string);(PVar "_17"%string);(PVar "_16"%string);(PVar "_15"%string);(PVar "_14"%string);(PVar "_13"%string);(PVar "_12"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_22"%string);(EVar "_21"%string);(EVar "_20"%string);(EVar "_19"%string);(EVar "_18"%string);(EVar "_17"%string);(EVar "_16"%string);(EVar "_15"%string);(EVar "_14"%string);(EVar "_13"%string);(EVar "_12"%string)])]))]) |};
          {| identifier := ("rukeymerge3_12b"%string, 12) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string;"_6"%string;"_7"%string;"_8"%string;"_9"%string;"_10"%string;"_11"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string);(EVar "_6"%string);(EVar "_7"%string);(EVar "_8"%string);(EVar "_9"%string);(EVar "_10"%string);(EVar "_11"%string)]) [([(PVar "I"%string);(PVar "E1"%string);(PVar "H1"%string);(PVar "T1"%string);(PVar "E2"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "E3"%string);(PVar "H3"%string);(PVar "T3"%string);(PVar "M"%string);(PVar "H2M"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "E2"%string);(EVar "E3"%string)]), (EApp (EFunId ("rukeymerge3_12_3"%string, 11)) [(EVar "I"%string);(EVar "E1"%string);(EVar "H1"%string);(EVar "T1"%string);(EVar "E2"%string);(EVar "H2"%string);(EVar "T2"%string);(ECons (EVar "H2M"%string) (EVar "M"%string));(EVar "E3"%string);(EVar "H3"%string);(EVar "T3"%string)]));([(PVar "I"%string);(PVar "E1"%string);(PVar "H1"%string);(PVar "T1"%string);(PVar "E2"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "E3"%string);(PVar "H3"%string);(PVar "T3"%string);(PVar "M"%string);(PVar "H2M"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rukeymerge3_2"%string, 11)) [(EVar "I"%string);(EVar "E1"%string);(EVar "H1"%string);(EVar "T1"%string);(EVar "T2"%string);(EVar "H2"%string);(EVar "E2"%string);(ECons (EVar "H2M"%string) (EVar "M"%string));(EVar "E3"%string);(EVar "H3"%string);(EVar "T3"%string)]))]) |};
          {| identifier := ("rukeymerge3_21b"%string, 12) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string;"_6"%string;"_7"%string;"_8"%string;"_9"%string;"_10"%string;"_11"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string);(EVar "_6"%string);(EVar "_7"%string);(EVar "_8"%string);(EVar "_9"%string);(EVar "_10"%string);(EVar "_11"%string)]) [([(PVar "I"%string);(PVar "E1"%string);(PVar "H1"%string);(PVar "T1"%string);(PVar "E2"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "E3"%string);(PVar "H3"%string);(PVar "T3"%string);(PVar "M"%string);(PVar "H2M"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "E1"%string);(EVar "E3"%string)]), (EApp (EFunId ("rukeymerge3_21_3"%string, 11)) [(EVar "I"%string);(EVar "E1"%string);(EVar "H1"%string);(EVar "T1"%string);(EVar "E2"%string);(EVar "H2"%string);(EVar "T2"%string);(ECons (EVar "H2M"%string) (EVar "M"%string));(EVar "E3"%string);(EVar "H3"%string);(EVar "T3"%string)]));([(PVar "I"%string);(PVar "_E1"%string);(PVar "H1"%string);(PVar "T1"%string);(PVar "E2"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "E3"%string);(PVar "H3"%string);(PVar "T3"%string);(PVar "M"%string);(PVar "H2M"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rukeymerge3_1"%string, 11)) [(EVar "I"%string);(EVar "T1"%string);(EVar "H1"%string);(EVar "T1"%string);(EVar "E2"%string);(EVar "H2"%string);(EVar "T2"%string);(ECons (EVar "H1"%string) (ECons (EVar "H2M"%string) (EVar "M"%string)));(EVar "E3"%string);(EVar "H3"%string);(EVar "T3"%string)]))]) |};
          {| identifier := ("rukeymerge3_12_3"%string, 11) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string;"_6"%string;"_7"%string;"_8"%string;"_9"%string;"_10"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string);(EVar "_6"%string);(EVar "_7"%string);(EVar "_8"%string);(EVar "_9"%string);(EVar "_10"%string)]) [([(PVar "I"%string);(PVar "E1"%string);(PVar "H1"%string);(PVar "T1"%string);(PVar "E2"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "M"%string);(PVar "E3M"%string);(PVar "H3M"%string);(PCons (PVar "H3"%string) (PVar "T3"%string))], (ELit (Atom "true"%string)), (ECase (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "I"%string);(EVar "H3"%string)]) [([(PVar "E3"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "E2"%string);(EVar "E3"%string)]), (EApp (EFunId ("rukeymerge3_12_3"%string, 11)) [(EVar "I"%string);(EVar "E1"%string);(EVar "H1"%string);(EVar "T1"%string);(EVar "E2"%string);(EVar "H2"%string);(EVar "T2"%string);(ECons (EVar "H3M"%string) (EVar "M"%string));(EVar "E3"%string);(EVar "H3"%string);(EVar "T3"%string)]));([(PVar "E3"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "E2"%string);(EVar "E3M"%string)]), (EApp (EFunId ("rukeymerge3_2"%string, 11)) [(EVar "I"%string);(EVar "E1"%string);(EVar "H1"%string);(EVar "T1"%string);(EVar "T2"%string);(EVar "H2"%string);(EVar "E2"%string);(EVar "M"%string);(EVar "E3"%string);(EVar "H3"%string);(EVar "T3"%string)]));([(PVar "E3"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rukeymerge3_2"%string, 11)) [(EVar "I"%string);(EVar "E1"%string);(EVar "H1"%string);(EVar "T1"%string);(EVar "T2"%string);(EVar "H2"%string);(EVar "E2"%string);(ECons (EVar "H3M"%string) (EVar "M"%string));(EVar "E3"%string);(EVar "H3"%string);(EVar "T3"%string)]))]));([(PVar "I"%string);(PVar "E1"%string);(PVar "H1"%string);(PVar "T1"%string);(PVar "E2"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "M"%string);(PVar "E3M"%string);(PVar "_H3M"%string);PNil], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "E2"%string);(EVar "E3M"%string)]), (EApp (EFunId ("rukeymerge2_2"%string, 8)) [(EVar "I"%string);(EVar "T1"%string);(EVar "E1"%string);(EVar "T2"%string);(EVar "M"%string);(EVar "E2"%string);(EVar "H2"%string);(EVar "H1"%string)]));([(PVar "I"%string);(PVar "E1"%string);(PVar "H1"%string);(PVar "T1"%string);(PVar "E2"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "M"%string);(PVar "_E3M"%string);(PVar "H3M"%string);PNil], (ELit (Atom "true"%string)), (EApp (EFunId ("rukeymerge2_2"%string, 8)) [(EVar "I"%string);(EVar "T1"%string);(EVar "E1"%string);(EVar "T2"%string);(ECons (EVar "H3M"%string) (EVar "M"%string));(EVar "E2"%string);(EVar "H2"%string);(EVar "H1"%string)]));([(PVar "_22"%string);(PVar "_21"%string);(PVar "_20"%string);(PVar "_19"%string);(PVar "_18"%string);(PVar "_17"%string);(PVar "_16"%string);(PVar "_15"%string);(PVar "_14"%string);(PVar "_13"%string);(PVar "_12"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_22"%string);(EVar "_21"%string);(EVar "_20"%string);(EVar "_19"%string);(EVar "_18"%string);(EVar "_17"%string);(EVar "_16"%string);(EVar "_15"%string);(EVar "_14"%string);(EVar "_13"%string);(EVar "_12"%string)])]))]) |};
          {| identifier := ("rukeymerge3_21_3"%string, 11) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string;"_6"%string;"_7"%string;"_8"%string;"_9"%string;"_10"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string);(EVar "_6"%string);(EVar "_7"%string);(EVar "_8"%string);(EVar "_9"%string);(EVar "_10"%string)]) [([(PVar "I"%string);(PVar "E1"%string);(PVar "H1"%string);(PVar "T1"%string);(PVar "E2"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "M"%string);(PVar "E3M"%string);(PVar "H3M"%string);(PCons (PVar "H3"%string) (PVar "T3"%string))], (ELit (Atom "true"%string)), (ECase (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "I"%string);(EVar "H3"%string)]) [([(PVar "E3"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "E1"%string);(EVar "E3"%string)]), (EApp (EFunId ("rukeymerge3_21_3"%string, 11)) [(EVar "I"%string);(EVar "E1"%string);(EVar "H1"%string);(EVar "T1"%string);(EVar "E2"%string);(EVar "H2"%string);(EVar "T2"%string);(ECons (EVar "H3M"%string) (EVar "M"%string));(EVar "E3"%string);(EVar "H3"%string);(EVar "T3"%string)]));([(PVar "E3"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "E1"%string);(EVar "E3M"%string)]), (EApp (EFunId ("rukeymerge3_1"%string, 11)) [(EVar "I"%string);(EVar "T1"%string);(EVar "H1"%string);(EVar "T1"%string);(EVar "E2"%string);(EVar "H2"%string);(EVar "T2"%string);(ECons (EVar "H1"%string) (EVar "M"%string));(EVar "E3"%string);(EVar "H3"%string);(EVar "T3"%string)]));([(PVar "E3"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rukeymerge3_1"%string, 11)) [(EVar "I"%string);(EVar "T1"%string);(EVar "H1"%string);(EVar "T1"%string);(EVar "E2"%string);(EVar "H2"%string);(EVar "T2"%string);(ECons (EVar "H1"%string) (ECons (EVar "H3M"%string) (EVar "M"%string)));(EVar "E3"%string);(EVar "H3"%string);(EVar "T3"%string)]))]));([(PVar "I"%string);(PVar "E1"%string);(PVar "H1"%string);(PVar "T1"%string);(PVar "E2"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "M"%string);(PVar "E3M"%string);(PVar "_H3M"%string);PNil], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "E1"%string);(EVar "E3M"%string)]), (EApp (EFunId ("rukeymerge2_1"%string, 6)) [(EVar "I"%string);(EVar "T1"%string);(EVar "E2"%string);(EVar "T2"%string);(ECons (EVar "H1"%string) (EVar "M"%string));(EVar "H2"%string)]));([(PVar "I"%string);(PVar "_E1"%string);(PVar "H1"%string);(PVar "T1"%string);(PVar "E2"%string);(PVar "H2"%string);(PVar "T2"%string);(PVar "M"%string);(PVar "_E3M"%string);(PVar "H3M"%string);PNil], (ELit (Atom "true"%string)), (EApp (EFunId ("rukeymerge2_1"%string, 6)) [(EVar "I"%string);(EVar "T1"%string);(EVar "E2"%string);(EVar "T2"%string);(ECons (EVar "H1"%string) (ECons (EVar "H3M"%string) (EVar "M"%string)));(EVar "H2"%string)]));([(PVar "_22"%string);(PVar "_21"%string);(PVar "_20"%string);(PVar "_19"%string);(PVar "_18"%string);(PVar "_17"%string);(PVar "_16"%string);(PVar "_15"%string);(PVar "_14"%string);(PVar "_13"%string);(PVar "_12"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_22"%string);(EVar "_21"%string);(EVar "_20"%string);(EVar "_19"%string);(EVar "_18"%string);(EVar "_17"%string);(EVar "_16"%string);(EVar "_15"%string);(EVar "_14"%string);(EVar "_13"%string);(EVar "_12"%string)])]))]) |};
          {| identifier := ("ukeymerge2_1"%string, 7) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string;"_6"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string);(EVar "_6"%string)]) [([(PVar "I"%string);(PCons (PVar "H1"%string) (PVar "T1"%string));(PVar "E2"%string);(PVar "HdM"%string);(PVar "T2"%string);(PVar "M"%string);(PVar "H2"%string)], (ELit (Atom "true"%string)), (ECase (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "I"%string);(EVar "H1"%string)]) [([(PVar "E1"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "E1"%string);(EVar "E2"%string)]), (EApp (EFunId ("ukeymerge2_1"%string, 7)) [(EVar "I"%string);(EVar "T1"%string);(EVar "E2"%string);(EVar "E1"%string);(EVar "T2"%string);(ECons (EVar "H1"%string) (EVar "M"%string));(EVar "H2"%string)]));([(PVar "E1"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "E2"%string);(EVar "HdM"%string)]), (EApp (EFunId ("ukeymerge2_2"%string, 6)) [(EVar "I"%string);(EVar "T1"%string);(EVar "E1"%string);(EVar "H1"%string);(EVar "T2"%string);(EVar "M"%string)]));([(PVar "E1"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("ukeymerge2_2"%string, 6)) [(EVar "I"%string);(EVar "T1"%string);(EVar "E1"%string);(EVar "H1"%string);(EVar "T2"%string);(ECons (EVar "H2"%string) (EVar "M"%string))]))]));([(PVar "_I"%string);PNil;(PVar "E2"%string);(PVar "HdM"%string);(PVar "T2"%string);(PVar "M"%string);(PVar "_H2"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "E2"%string);(EVar "HdM"%string)]), (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "T2"%string);(EVar "M"%string)]));([(PVar "_I"%string);PNil;(PVar "_E2"%string);(PVar "_HdM"%string);(PVar "T2"%string);(PVar "M"%string);(PVar "H2"%string)], (ELit (Atom "true"%string)), (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "T2"%string);(ECons (EVar "H2"%string) (EVar "M"%string))]));([(PVar "_14"%string);(PVar "_13"%string);(PVar "_12"%string);(PVar "_11"%string);(PVar "_10"%string);(PVar "_9"%string);(PVar "_8"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_14"%string);(EVar "_13"%string);(EVar "_12"%string);(EVar "_11"%string);(EVar "_10"%string);(EVar "_9"%string);(EVar "_8"%string)])]))]) |};
          {| identifier := ("ukeymerge2_2"%string, 6) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string)]) [([(PVar "I"%string);(PVar "T1"%string);(PVar "E1"%string);(PVar "H1"%string);(PCons (PVar "H2"%string) (PVar "T2"%string));(PVar "M"%string)], (ELit (Atom "true"%string)), (ECase (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "I"%string);(EVar "H2"%string)]) [([(PVar "E2"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "E1"%string);(EVar "E2"%string)]), (EApp (EFunId ("ukeymerge2_1"%string, 7)) [(EVar "I"%string);(EVar "T1"%string);(EVar "E2"%string);(EVar "E1"%string);(EVar "T2"%string);(ECons (EVar "H1"%string) (EVar "M"%string));(EVar "H2"%string)]));([(PVar "_E2"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("ukeymerge2_2"%string, 6)) [(EVar "I"%string);(EVar "T1"%string);(EVar "E1"%string);(EVar "H1"%string);(EVar "T2"%string);(ECons (EVar "H2"%string) (EVar "M"%string))]))]));([(PVar "_I"%string);(PVar "T1"%string);(PVar "_E1"%string);(PVar "H1"%string);PNil;(PVar "M"%string)], (ELit (Atom "true"%string)), (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "T1"%string);(ECons (EVar "H1"%string) (EVar "M"%string))]));([(PVar "_12"%string);(PVar "_11"%string);(PVar "_10"%string);(PVar "_9"%string);(PVar "_8"%string);(PVar "_7"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_12"%string);(EVar "_11"%string);(EVar "_10"%string);(EVar "_9"%string);(EVar "_8"%string);(EVar "_7"%string)])]))]) |};
          {| identifier := ("rukeymerge2_1"%string, 6) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string)]) [([(PVar "I"%string);(PCons (PVar "H1"%string) (PVar "T1"%string));(PVar "E2"%string);(PVar "T2"%string);(PVar "M"%string);(PVar "H2"%string)], (ELit (Atom "true"%string)), (ECase (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "I"%string);(EVar "H1"%string)]) [([(PVar "E1"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "E1"%string);(EVar "E2"%string)]), (EApp (EFunId ("rukeymerge2_2"%string, 8)) [(EVar "I"%string);(EVar "T1"%string);(EVar "E1"%string);(EVar "T2"%string);(EVar "M"%string);(EVar "E2"%string);(EVar "H2"%string);(EVar "H1"%string)]));([(PVar "_E1"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rukeymerge2_1"%string, 6)) [(EVar "I"%string);(EVar "T1"%string);(EVar "E2"%string);(EVar "T2"%string);(ECons (EVar "H1"%string) (EVar "M"%string));(EVar "H2"%string)]))]));([(PVar "_I"%string);PNil;(PVar "_E2"%string);(PVar "T2"%string);(PVar "M"%string);(PVar "H2"%string)], (ELit (Atom "true"%string)), (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "T2"%string);(ECons (EVar "H2"%string) (EVar "M"%string))]));([(PVar "_12"%string);(PVar "_11"%string);(PVar "_10"%string);(PVar "_9"%string);(PVar "_8"%string);(PVar "_7"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_12"%string);(EVar "_11"%string);(EVar "_10"%string);(EVar "_9"%string);(EVar "_8"%string);(EVar "_7"%string)])]))]) |};
          {| identifier := ("rukeymerge2_2"%string, 8) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string;"_6"%string;"_7"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string);(EVar "_6"%string);(EVar "_7"%string)]) [([(PVar "I"%string);(PVar "T1"%string);(PVar "E1"%string);(PCons (PVar "H2"%string) (PVar "T2"%string));(PVar "M"%string);(PVar "E2M"%string);(PVar "H2M"%string);(PVar "H1"%string)], (ELit (Atom "true"%string)), (ECase (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "element"%string)) [(EVar "I"%string);(EVar "H2"%string)]) [([(PVar "E2"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=<"%string)) [(EVar "E1"%string);(EVar "E2"%string)]), (EApp (EFunId ("rukeymerge2_2"%string, 8)) [(EVar "I"%string);(EVar "T1"%string);(EVar "E1"%string);(EVar "T2"%string);(ECons (EVar "H2M"%string) (EVar "M"%string));(EVar "E2"%string);(EVar "H2"%string);(EVar "H1"%string)]));([(PVar "E2"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "E1"%string);(EVar "E2M"%string)]), (EApp (EFunId ("rukeymerge2_1"%string, 6)) [(EVar "I"%string);(EVar "T1"%string);(EVar "E2"%string);(EVar "T2"%string);(ECons (EVar "H1"%string) (EVar "M"%string));(EVar "H2"%string)]));([(PVar "E2"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rukeymerge2_1"%string, 6)) [(EVar "I"%string);(EVar "T1"%string);(EVar "E2"%string);(EVar "T2"%string);(ECons (EVar "H1"%string) (ECons (EVar "H2M"%string) (EVar "M"%string)));(EVar "H2"%string)]))]));([(PVar "_I"%string);(PVar "T1"%string);(PVar "E1"%string);PNil;(PVar "M"%string);(PVar "E2M"%string);(PVar "_H2M"%string);(PVar "H1"%string)], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "E1"%string);(EVar "E2M"%string)]), (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "T1"%string);(ECons (EVar "H1"%string) (EVar "M"%string))]));([(PVar "_I"%string);(PVar "T1"%string);(PVar "_E1"%string);PNil;(PVar "M"%string);(PVar "_E2M"%string);(PVar "H2M"%string);(PVar "H1"%string)], (ELit (Atom "true"%string)), (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "T1"%string);(ECons (EVar "H1"%string) (ECons (EVar "H2M"%string) (EVar "M"%string)))]));([(PVar "_16"%string);(PVar "_15"%string);(PVar "_14"%string);(PVar "_13"%string);(PVar "_12"%string);(PVar "_11"%string);(PVar "_10"%string);(PVar "_9"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_16"%string);(EVar "_15"%string);(EVar "_14"%string);(EVar "_13"%string);(EVar "_12"%string);(EVar "_11"%string);(EVar "_10"%string);(EVar "_9"%string)])]))]) |};
          {| identifier := ("fsplit_1"%string, 6) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string)]) [([(PVar "Y"%string);(PVar "X"%string);(PVar "Fun"%string);(PCons (PVar "Z"%string) (PVar "L"%string));(PVar "R"%string);(PVar "Rs"%string)], (ELit (Atom "true"%string)), (ECase (EApp (EVar "Fun"%string) [(EVar "Y"%string);(EVar "Z"%string)]) [([(PLit (Atom "true"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("fsplit_1"%string, 6)) [(EVar "Z"%string);(EVar "Y"%string);(EVar "Fun"%string);(EVar "L"%string);(ECons (EVar "X"%string) (EVar "R"%string));(EVar "Rs"%string)]));([(PLit (Atom "false"%string))], (ELit (Atom "true"%string)), (ECase (EApp (EVar "Fun"%string) [(EVar "X"%string);(EVar "Z"%string)]) [([(PLit (Atom "true"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("fsplit_1"%string, 6)) [(EVar "Y"%string);(EVar "Z"%string);(EVar "Fun"%string);(EVar "L"%string);(ECons (EVar "X"%string) (EVar "R"%string));(EVar "Rs"%string)]));([(PLit (Atom "false"%string))], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "R"%string);ENil]), (EApp (EFunId ("fsplit_1"%string, 6)) [(EVar "Y"%string);(EVar "X"%string);(EVar "Fun"%string);(EVar "L"%string);(ECons (EVar "Z"%string) ENil);(EVar "Rs"%string)]));([(PLit (Atom "false"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("fsplit_1_1"%string, 7)) [(EVar "Y"%string);(EVar "X"%string);(EVar "Fun"%string);(EVar "L"%string);(EVar "R"%string);(EVar "Rs"%string);(EVar "Z"%string)]));([(PVar "_6"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "case_clause"%string));(EVar "_6"%string)])]))]));([(PVar "_7"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "case_clause"%string));(EVar "_7"%string)])]))]));([(PVar "Y"%string);(PVar "X"%string);(PVar "Fun"%string);PNil;(PVar "R"%string);(PVar "Rs"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rfmergel"%string, 4)) [(ECons (ECons (EVar "Y"%string) (ECons (EVar "X"%string) (EVar "R"%string))) (EVar "Rs"%string));ENil;(EVar "Fun"%string);(ELit (Atom "asc"%string))]));([(PVar "_13"%string);(PVar "_12"%string);(PVar "_11"%string);(PVar "_10"%string);(PVar "_9"%string);(PVar "_8"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_13"%string);(EVar "_12"%string);(EVar "_11"%string);(EVar "_10"%string);(EVar "_9"%string);(EVar "_8"%string)])]))]) |};
          {| identifier := ("fsplit_1_1"%string, 7) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string;"_6"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string);(EVar "_6"%string)]) [([(PVar "Y"%string);(PVar "X"%string);(PVar "Fun"%string);(PCons (PVar "Z"%string) (PVar "L"%string));(PVar "R"%string);(PVar "Rs"%string);(PVar "S"%string)], (ELit (Atom "true"%string)), (ECase (EApp (EVar "Fun"%string) [(EVar "Y"%string);(EVar "Z"%string)]) [([(PLit (Atom "true"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("fsplit_1_1"%string, 7)) [(EVar "Z"%string);(EVar "Y"%string);(EVar "Fun"%string);(EVar "L"%string);(ECons (EVar "X"%string) (EVar "R"%string));(EVar "Rs"%string);(EVar "S"%string)]));([(PLit (Atom "false"%string))], (ELit (Atom "true"%string)), (ECase (EApp (EVar "Fun"%string) [(EVar "X"%string);(EVar "Z"%string)]) [([(PLit (Atom "true"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("fsplit_1_1"%string, 7)) [(EVar "Y"%string);(EVar "Z"%string);(EVar "Fun"%string);(EVar "L"%string);(ECons (EVar "X"%string) (EVar "R"%string));(EVar "Rs"%string);(EVar "S"%string)]));([(PLit (Atom "false"%string))], (ELit (Atom "true"%string)), (ECase (EApp (EVar "Fun"%string) [(EVar "S"%string);(EVar "Z"%string)]) [([(PLit (Atom "true"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("fsplit_1"%string, 6)) [(EVar "Z"%string);(EVar "S"%string);(EVar "Fun"%string);(EVar "L"%string);ENil;(ECons (ECons (EVar "Y"%string) (ECons (EVar "X"%string) (EVar "R"%string))) (EVar "Rs"%string))]));([(PLit (Atom "false"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("fsplit_1"%string, 6)) [(EVar "S"%string);(EVar "Z"%string);(EVar "Fun"%string);(EVar "L"%string);ENil;(ECons (ECons (EVar "Y"%string) (ECons (EVar "X"%string) (EVar "R"%string))) (EVar "Rs"%string))]));([(PVar "_7"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "case_clause"%string));(EVar "_7"%string)])]))]));([(PVar "_8"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "case_clause"%string));(EVar "_8"%string)])]))]));([(PVar "_9"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "case_clause"%string));(EVar "_9"%string)])]))]));([(PVar "Y"%string);(PVar "X"%string);(PVar "Fun"%string);PNil;(PVar "R"%string);(PVar "Rs"%string);(PVar "S"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rfmergel"%string, 4)) [(ECons (ECons (EVar "S"%string) ENil) (ECons (ECons (EVar "Y"%string) (ECons (EVar "X"%string) (EVar "R"%string))) (EVar "Rs"%string)));ENil;(EVar "Fun"%string);(ELit (Atom "asc"%string))]));([(PVar "_16"%string);(PVar "_15"%string);(PVar "_14"%string);(PVar "_13"%string);(PVar "_12"%string);(PVar "_11"%string);(PVar "_10"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_16"%string);(EVar "_15"%string);(EVar "_14"%string);(EVar "_13"%string);(EVar "_12"%string);(EVar "_11"%string);(EVar "_10"%string)])]))]) |};
          {| identifier := ("fsplit_2"%string, 6) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string)]) [([(PVar "Y"%string);(PVar "X"%string);(PVar "Fun"%string);(PCons (PVar "Z"%string) (PVar "L"%string));(PVar "R"%string);(PVar "Rs"%string)], (ELit (Atom "true"%string)), (ECase (EApp (EVar "Fun"%string) [(EVar "Y"%string);(EVar "Z"%string)]) [([(PLit (Atom "false"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("fsplit_2"%string, 6)) [(EVar "Z"%string);(EVar "Y"%string);(EVar "Fun"%string);(EVar "L"%string);(ECons (EVar "X"%string) (EVar "R"%string));(EVar "Rs"%string)]));([(PLit (Atom "true"%string))], (ELit (Atom "true"%string)), (ECase (EApp (EVar "Fun"%string) [(EVar "X"%string);(EVar "Z"%string)]) [([(PLit (Atom "false"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("fsplit_2"%string, 6)) [(EVar "Y"%string);(EVar "Z"%string);(EVar "Fun"%string);(EVar "L"%string);(ECons (EVar "X"%string) (EVar "R"%string));(EVar "Rs"%string)]));([(PLit (Atom "true"%string))], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "R"%string);ENil]), (EApp (EFunId ("fsplit_2"%string, 6)) [(EVar "Y"%string);(EVar "X"%string);(EVar "Fun"%string);(EVar "L"%string);(ECons (EVar "Z"%string) ENil);(EVar "Rs"%string)]));([(PLit (Atom "true"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("fsplit_2_1"%string, 7)) [(EVar "Y"%string);(EVar "X"%string);(EVar "Fun"%string);(EVar "L"%string);(EVar "R"%string);(EVar "Rs"%string);(EVar "Z"%string)]));([(PVar "_6"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "case_clause"%string));(EVar "_6"%string)])]))]));([(PVar "_7"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "case_clause"%string));(EVar "_7"%string)])]))]));([(PVar "Y"%string);(PVar "X"%string);(PVar "Fun"%string);PNil;(PVar "R"%string);(PVar "Rs"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("fmergel"%string, 4)) [(ECons (ECons (EVar "Y"%string) (ECons (EVar "X"%string) (EVar "R"%string))) (EVar "Rs"%string));ENil;(EVar "Fun"%string);(ELit (Atom "desc"%string))]));([(PVar "_13"%string);(PVar "_12"%string);(PVar "_11"%string);(PVar "_10"%string);(PVar "_9"%string);(PVar "_8"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_13"%string);(EVar "_12"%string);(EVar "_11"%string);(EVar "_10"%string);(EVar "_9"%string);(EVar "_8"%string)])]))]) |};
          {| identifier := ("fsplit_2_1"%string, 7) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string;"_6"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string);(EVar "_6"%string)]) [([(PVar "Y"%string);(PVar "X"%string);(PVar "Fun"%string);(PCons (PVar "Z"%string) (PVar "L"%string));(PVar "R"%string);(PVar "Rs"%string);(PVar "S"%string)], (ELit (Atom "true"%string)), (ECase (EApp (EVar "Fun"%string) [(EVar "Y"%string);(EVar "Z"%string)]) [([(PLit (Atom "false"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("fsplit_2_1"%string, 7)) [(EVar "Z"%string);(EVar "Y"%string);(EVar "Fun"%string);(EVar "L"%string);(ECons (EVar "X"%string) (EVar "R"%string));(EVar "Rs"%string);(EVar "S"%string)]));([(PLit (Atom "true"%string))], (ELit (Atom "true"%string)), (ECase (EApp (EVar "Fun"%string) [(EVar "X"%string);(EVar "Z"%string)]) [([(PLit (Atom "false"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("fsplit_2_1"%string, 7)) [(EVar "Y"%string);(EVar "Z"%string);(EVar "Fun"%string);(EVar "L"%string);(ECons (EVar "X"%string) (EVar "R"%string));(EVar "Rs"%string);(EVar "S"%string)]));([(PLit (Atom "true"%string))], (ELit (Atom "true"%string)), (ECase (EApp (EVar "Fun"%string) [(EVar "S"%string);(EVar "Z"%string)]) [([(PLit (Atom "false"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("fsplit_2"%string, 6)) [(EVar "Z"%string);(EVar "S"%string);(EVar "Fun"%string);(EVar "L"%string);ENil;(ECons (ECons (EVar "Y"%string) (ECons (EVar "X"%string) (EVar "R"%string))) (EVar "Rs"%string))]));([(PLit (Atom "true"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("fsplit_2"%string, 6)) [(EVar "S"%string);(EVar "Z"%string);(EVar "Fun"%string);(EVar "L"%string);ENil;(ECons (ECons (EVar "Y"%string) (ECons (EVar "X"%string) (EVar "R"%string))) (EVar "Rs"%string))]));([(PVar "_7"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "case_clause"%string));(EVar "_7"%string)])]))]));([(PVar "_8"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "case_clause"%string));(EVar "_8"%string)])]))]));([(PVar "_9"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "case_clause"%string));(EVar "_9"%string)])]))]));([(PVar "Y"%string);(PVar "X"%string);(PVar "Fun"%string);PNil;(PVar "R"%string);(PVar "Rs"%string);(PVar "S"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("fmergel"%string, 4)) [(ECons (ECons (EVar "S"%string) ENil) (ECons (ECons (EVar "Y"%string) (ECons (EVar "X"%string) (EVar "R"%string))) (EVar "Rs"%string)));ENil;(EVar "Fun"%string);(ELit (Atom "desc"%string))]));([(PVar "_16"%string);(PVar "_15"%string);(PVar "_14"%string);(PVar "_13"%string);(PVar "_12"%string);(PVar "_11"%string);(PVar "_10"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_16"%string);(EVar "_15"%string);(EVar "_14"%string);(EVar "_13"%string);(EVar "_12"%string);(EVar "_11"%string);(EVar "_10"%string)])]))]) |};
          {| identifier := ("fmergel"%string, 4) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string)]) [([(PCons (PVar "T1"%string) (PCons (PCons (PVar "H2"%string) (PVar "T2"%string)) (PVar "L"%string)));(PVar "Acc"%string);(PVar "Fun"%string);(PLit (Atom "asc"%string))], (ELit (Atom "true"%string)), (ELet ["_4"%string] (EApp (EFunId ("fmerge2_1"%string, 5)) [(EVar "T1"%string);(EVar "H2"%string);(EVar "Fun"%string);(EVar "T2"%string);ENil]) (EApp (EFunId ("fmergel"%string, 4)) [(EVar "L"%string);(ECons (EVar "_4"%string) (EVar "Acc"%string));(EVar "Fun"%string);(ELit (Atom "asc"%string))])));([(PCons (PCons (PVar "H2"%string) (PVar "T2"%string)) (PCons (PVar "T1"%string) (PVar "L"%string)));(PVar "Acc"%string);(PVar "Fun"%string);(PLit (Atom "desc"%string))], (ELit (Atom "true"%string)), (ELet ["_5"%string] (EApp (EFunId ("fmerge2_1"%string, 5)) [(EVar "T1"%string);(EVar "H2"%string);(EVar "Fun"%string);(EVar "T2"%string);ENil]) (EApp (EFunId ("fmergel"%string, 4)) [(EVar "L"%string);(ECons (EVar "_5"%string) (EVar "Acc"%string));(EVar "Fun"%string);(ELit (Atom "desc"%string))])));([(PCons (PVar "L"%string) PNil);PNil;(PVar "_Fun"%string);(PVar "_O"%string)], (ELit (Atom "true"%string)), (EVar "L"%string));([(PCons (PVar "L"%string) PNil);(PVar "Acc"%string);(PVar "Fun"%string);(PVar "O"%string)], (ELit (Atom "true"%string)), (ELet ["_6"%string] (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "L"%string);ENil]) (EApp (EFunId ("rfmergel"%string, 4)) [(ECons (EVar "_6"%string) (EVar "Acc"%string));ENil;(EVar "Fun"%string);(EVar "O"%string)])));([PNil;(PVar "Acc"%string);(PVar "Fun"%string);(PVar "O"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rfmergel"%string, 4)) [(EVar "Acc"%string);ENil;(EVar "Fun"%string);(EVar "O"%string)]));([(PVar "_10"%string);(PVar "_9"%string);(PVar "_8"%string);(PVar "_7"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_10"%string);(EVar "_9"%string);(EVar "_8"%string);(EVar "_7"%string)])]))]) |};
          {| identifier := ("rfmergel"%string, 4) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string)]) [([(PCons (PCons (PVar "H2"%string) (PVar "T2"%string)) (PCons (PVar "T1"%string) (PVar "L"%string)));(PVar "Acc"%string);(PVar "Fun"%string);(PLit (Atom "asc"%string))], (ELit (Atom "true"%string)), (ELet ["_4"%string] (EApp (EFunId ("rfmerge2_1"%string, 5)) [(EVar "T1"%string);(EVar "H2"%string);(EVar "Fun"%string);(EVar "T2"%string);ENil]) (EApp (EFunId ("rfmergel"%string, 4)) [(EVar "L"%string);(ECons (EVar "_4"%string) (EVar "Acc"%string));(EVar "Fun"%string);(ELit (Atom "asc"%string))])));([(PCons (PVar "T1"%string) (PCons (PCons (PVar "H2"%string) (PVar "T2"%string)) (PVar "L"%string)));(PVar "Acc"%string);(PVar "Fun"%string);(PLit (Atom "desc"%string))], (ELit (Atom "true"%string)), (ELet ["_5"%string] (EApp (EFunId ("rfmerge2_1"%string, 5)) [(EVar "T1"%string);(EVar "H2"%string);(EVar "Fun"%string);(EVar "T2"%string);ENil]) (EApp (EFunId ("rfmergel"%string, 4)) [(EVar "L"%string);(ECons (EVar "_5"%string) (EVar "Acc"%string));(EVar "Fun"%string);(ELit (Atom "desc"%string))])));([(PCons (PVar "L"%string) PNil);(PVar "Acc"%string);(PVar "Fun"%string);(PVar "O"%string)], (ELit (Atom "true"%string)), (ELet ["_6"%string] (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "L"%string);ENil]) (EApp (EFunId ("fmergel"%string, 4)) [(ECons (EVar "_6"%string) (EVar "Acc"%string));ENil;(EVar "Fun"%string);(EVar "O"%string)])));([PNil;(PVar "Acc"%string);(PVar "Fun"%string);(PVar "O"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("fmergel"%string, 4)) [(EVar "Acc"%string);ENil;(EVar "Fun"%string);(EVar "O"%string)]));([(PVar "_10"%string);(PVar "_9"%string);(PVar "_8"%string);(PVar "_7"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_10"%string);(EVar "_9"%string);(EVar "_8"%string);(EVar "_7"%string)])]))]) |};
          {| identifier := ("fmerge2_1"%string, 5) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string)]) [([(PCons (PVar "H1"%string) (PVar "T1"%string));(PVar "H2"%string);(PVar "Fun"%string);(PVar "T2"%string);(PVar "M"%string)], (ELit (Atom "true"%string)), (ECase (EApp (EVar "Fun"%string) [(EVar "H1"%string);(EVar "H2"%string)]) [([(PLit (Atom "true"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("fmerge2_1"%string, 5)) [(EVar "T1"%string);(EVar "H2"%string);(EVar "Fun"%string);(EVar "T2"%string);(ECons (EVar "H1"%string) (EVar "M"%string))]));([(PLit (Atom "false"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("fmerge2_2"%string, 5)) [(EVar "H1"%string);(EVar "T1"%string);(EVar "Fun"%string);(EVar "T2"%string);(ECons (EVar "H2"%string) (EVar "M"%string))]));([(PVar "_5"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "case_clause"%string));(EVar "_5"%string)])]))]));([PNil;(PVar "H2"%string);(PVar "_Fun"%string);(PVar "T2"%string);(PVar "M"%string)], (ELit (Atom "true"%string)), (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "T2"%string);(ECons (EVar "H2"%string) (EVar "M"%string))]));([(PVar "_10"%string);(PVar "_9"%string);(PVar "_8"%string);(PVar "_7"%string);(PVar "_6"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_10"%string);(EVar "_9"%string);(EVar "_8"%string);(EVar "_7"%string);(EVar "_6"%string)])]))]) |};
          {| identifier := ("fmerge2_2"%string, 5) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string)]) [([(PVar "H1"%string);(PVar "T1"%string);(PVar "Fun"%string);(PCons (PVar "H2"%string) (PVar "T2"%string));(PVar "M"%string)], (ELit (Atom "true"%string)), (ECase (EApp (EVar "Fun"%string) [(EVar "H1"%string);(EVar "H2"%string)]) [([(PLit (Atom "true"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("fmerge2_1"%string, 5)) [(EVar "T1"%string);(EVar "H2"%string);(EVar "Fun"%string);(EVar "T2"%string);(ECons (EVar "H1"%string) (EVar "M"%string))]));([(PLit (Atom "false"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("fmerge2_2"%string, 5)) [(EVar "H1"%string);(EVar "T1"%string);(EVar "Fun"%string);(EVar "T2"%string);(ECons (EVar "H2"%string) (EVar "M"%string))]));([(PVar "_5"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "case_clause"%string));(EVar "_5"%string)])]))]));([(PVar "H1"%string);(PVar "T1"%string);(PVar "_Fun"%string);PNil;(PVar "M"%string)], (ELit (Atom "true"%string)), (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "T1"%string);(ECons (EVar "H1"%string) (EVar "M"%string))]));([(PVar "_10"%string);(PVar "_9"%string);(PVar "_8"%string);(PVar "_7"%string);(PVar "_6"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_10"%string);(EVar "_9"%string);(EVar "_8"%string);(EVar "_7"%string);(EVar "_6"%string)])]))]) |};
          {| identifier := ("rfmerge2_1"%string, 5) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string)]) [([(PCons (PVar "H1"%string) (PVar "T1"%string));(PVar "H2"%string);(PVar "Fun"%string);(PVar "T2"%string);(PVar "M"%string)], (ELit (Atom "true"%string)), (ECase (EApp (EVar "Fun"%string) [(EVar "H1"%string);(EVar "H2"%string)]) [([(PLit (Atom "true"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("rfmerge2_2"%string, 5)) [(EVar "H1"%string);(EVar "T1"%string);(EVar "Fun"%string);(EVar "T2"%string);(ECons (EVar "H2"%string) (EVar "M"%string))]));([(PLit (Atom "false"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("rfmerge2_1"%string, 5)) [(EVar "T1"%string);(EVar "H2"%string);(EVar "Fun"%string);(EVar "T2"%string);(ECons (EVar "H1"%string) (EVar "M"%string))]));([(PVar "_5"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "case_clause"%string));(EVar "_5"%string)])]))]));([PNil;(PVar "H2"%string);(PVar "_Fun"%string);(PVar "T2"%string);(PVar "M"%string)], (ELit (Atom "true"%string)), (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "T2"%string);(ECons (EVar "H2"%string) (EVar "M"%string))]));([(PVar "_10"%string);(PVar "_9"%string);(PVar "_8"%string);(PVar "_7"%string);(PVar "_6"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_10"%string);(EVar "_9"%string);(EVar "_8"%string);(EVar "_7"%string);(EVar "_6"%string)])]))]) |};
          {| identifier := ("rfmerge2_2"%string, 5) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string)]) [([(PVar "H1"%string);(PVar "T1"%string);(PVar "Fun"%string);(PCons (PVar "H2"%string) (PVar "T2"%string));(PVar "M"%string)], (ELit (Atom "true"%string)), (ECase (EApp (EVar "Fun"%string) [(EVar "H1"%string);(EVar "H2"%string)]) [([(PLit (Atom "true"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("rfmerge2_2"%string, 5)) [(EVar "H1"%string);(EVar "T1"%string);(EVar "Fun"%string);(EVar "T2"%string);(ECons (EVar "H2"%string) (EVar "M"%string))]));([(PLit (Atom "false"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("rfmerge2_1"%string, 5)) [(EVar "T1"%string);(EVar "H2"%string);(EVar "Fun"%string);(EVar "T2"%string);(ECons (EVar "H1"%string) (EVar "M"%string))]));([(PVar "_5"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "case_clause"%string));(EVar "_5"%string)])]))]));([(PVar "H1"%string);(PVar "T1"%string);(PVar "_Fun"%string);PNil;(PVar "M"%string)], (ELit (Atom "true"%string)), (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "T1"%string);(ECons (EVar "H1"%string) (EVar "M"%string))]));([(PVar "_10"%string);(PVar "_9"%string);(PVar "_8"%string);(PVar "_7"%string);(PVar "_6"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_10"%string);(EVar "_9"%string);(EVar "_8"%string);(EVar "_7"%string);(EVar "_6"%string)])]))]) |};
          {| identifier := ("ufsplit_1"%string, 6) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string)]) [([(PVar "Y"%string);(PVar "X"%string);(PVar "Fun"%string);(PCons (PVar "Z"%string) (PVar "L"%string));(PVar "R"%string);(PVar "Rs"%string)], (ELit (Atom "true"%string)), (ECase (EApp (EVar "Fun"%string) [(EVar "Y"%string);(EVar "Z"%string)]) [([(PLit (Atom "true"%string))], (ELit (Atom "true"%string)), (ECase (EApp (EVar "Fun"%string) [(EVar "Z"%string);(EVar "Y"%string)]) [([(PLit (Atom "true"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("ufsplit_1"%string, 6)) [(EVar "Y"%string);(EVar "X"%string);(EVar "Fun"%string);(EVar "L"%string);(EVar "R"%string);(EVar "Rs"%string)]));([(PLit (Atom "false"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("ufsplit_1"%string, 6)) [(EVar "Z"%string);(EVar "Y"%string);(EVar "Fun"%string);(EVar "L"%string);(ECons (EVar "X"%string) (EVar "R"%string));(EVar "Rs"%string)]));([(PVar "_6"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "case_clause"%string));(EVar "_6"%string)])]))]));([(PLit (Atom "false"%string))], (ELit (Atom "true"%string)), (ECase (EApp (EVar "Fun"%string) [(EVar "X"%string);(EVar "Z"%string)]) [([(PLit (Atom "true"%string))], (ELit (Atom "true"%string)), (ECase (EApp (EVar "Fun"%string) [(EVar "Z"%string);(EVar "X"%string)]) [([(PLit (Atom "true"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("ufsplit_1"%string, 6)) [(EVar "Y"%string);(EVar "X"%string);(EVar "Fun"%string);(EVar "L"%string);(EVar "R"%string);(EVar "Rs"%string)]));([(PLit (Atom "false"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("ufsplit_1"%string, 6)) [(EVar "Y"%string);(EVar "Z"%string);(EVar "Fun"%string);(EVar "L"%string);(ECons (EVar "X"%string) (EVar "R"%string));(EVar "Rs"%string)]));([(PVar "_7"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "case_clause"%string));(EVar "_7"%string)])]))]));([(PLit (Atom "false"%string))], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=="%string)) [(EVar "R"%string);ENil]), (EApp (EFunId ("ufsplit_1"%string, 6)) [(EVar "Y"%string);(EVar "X"%string);(EVar "Fun"%string);(EVar "L"%string);(ECons (EVar "Z"%string) ENil);(EVar "Rs"%string)]));([(PLit (Atom "false"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("ufsplit_1_1"%string, 7)) [(EVar "Y"%string);(EVar "X"%string);(EVar "Fun"%string);(EVar "L"%string);(EVar "R"%string);(EVar "Rs"%string);(EVar "Z"%string)]));([(PVar "_8"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "case_clause"%string));(EVar "_8"%string)])]))]));([(PVar "_9"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "case_clause"%string));(EVar "_9"%string)])]))]));([(PVar "Y"%string);(PVar "X"%string);(PVar "Fun"%string);PNil;(PVar "R"%string);(PVar "Rs"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rufmergel"%string, 3)) [(ECons (ECons (EVar "Y"%string) (ECons (EVar "X"%string) (EVar "R"%string))) (EVar "Rs"%string));ENil;(EVar "Fun"%string)]));([(PVar "_15"%string);(PVar "_14"%string);(PVar "_13"%string);(PVar "_12"%string);(PVar "_11"%string);(PVar "_10"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_15"%string);(EVar "_14"%string);(EVar "_13"%string);(EVar "_12"%string);(EVar "_11"%string);(EVar "_10"%string)])]))]) |};
          {| identifier := ("ufsplit_1_1"%string, 7) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string;"_6"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string);(EVar "_6"%string)]) [([(PVar "Y"%string);(PVar "X"%string);(PVar "Fun"%string);(PCons (PVar "Z"%string) (PVar "L"%string));(PVar "R"%string);(PVar "Rs"%string);(PVar "S"%string)], (ELit (Atom "true"%string)), (ECase (EApp (EVar "Fun"%string) [(EVar "Y"%string);(EVar "Z"%string)]) [([(PLit (Atom "true"%string))], (ELit (Atom "true"%string)), (ECase (EApp (EVar "Fun"%string) [(EVar "Z"%string);(EVar "Y"%string)]) [([(PLit (Atom "true"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("ufsplit_1_1"%string, 7)) [(EVar "Y"%string);(EVar "X"%string);(EVar "Fun"%string);(EVar "L"%string);(EVar "R"%string);(EVar "Rs"%string);(EVar "S"%string)]));([(PLit (Atom "false"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("ufsplit_1_1"%string, 7)) [(EVar "Z"%string);(EVar "Y"%string);(EVar "Fun"%string);(EVar "L"%string);(ECons (EVar "X"%string) (EVar "R"%string));(EVar "Rs"%string);(EVar "S"%string)]));([(PVar "_7"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "case_clause"%string));(EVar "_7"%string)])]))]));([(PLit (Atom "false"%string))], (ELit (Atom "true"%string)), (ECase (EApp (EVar "Fun"%string) [(EVar "X"%string);(EVar "Z"%string)]) [([(PLit (Atom "true"%string))], (ELit (Atom "true"%string)), (ECase (EApp (EVar "Fun"%string) [(EVar "Z"%string);(EVar "X"%string)]) [([(PLit (Atom "true"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("ufsplit_1_1"%string, 7)) [(EVar "Y"%string);(EVar "X"%string);(EVar "Fun"%string);(EVar "L"%string);(EVar "R"%string);(EVar "Rs"%string);(EVar "S"%string)]));([(PLit (Atom "false"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("ufsplit_1_1"%string, 7)) [(EVar "Y"%string);(EVar "Z"%string);(EVar "Fun"%string);(EVar "L"%string);(ECons (EVar "X"%string) (EVar "R"%string));(EVar "Rs"%string);(EVar "S"%string)]));([(PVar "_8"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "case_clause"%string));(EVar "_8"%string)])]))]));([(PLit (Atom "false"%string))], (ELit (Atom "true"%string)), (ECase (EApp (EVar "Fun"%string) [(EVar "S"%string);(EVar "Z"%string)]) [([(PLit (Atom "true"%string))], (ELit (Atom "true"%string)), (ECase (EApp (EVar "Fun"%string) [(EVar "Z"%string);(EVar "S"%string)]) [([(PLit (Atom "true"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("ufsplit_1_1"%string, 7)) [(EVar "Y"%string);(EVar "X"%string);(EVar "Fun"%string);(EVar "L"%string);(EVar "R"%string);(EVar "Rs"%string);(EVar "S"%string)]));([(PLit (Atom "false"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("ufsplit_1"%string, 6)) [(EVar "Z"%string);(EVar "S"%string);(EVar "Fun"%string);(EVar "L"%string);ENil;(ECons (ECons (EVar "Y"%string) (ECons (EVar "X"%string) (EVar "R"%string))) (EVar "Rs"%string))]));([(PVar "_9"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "case_clause"%string));(EVar "_9"%string)])]))]));([(PLit (Atom "false"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("ufsplit_1"%string, 6)) [(EVar "S"%string);(EVar "Z"%string);(EVar "Fun"%string);(EVar "L"%string);ENil;(ECons (ECons (EVar "Y"%string) (ECons (EVar "X"%string) (EVar "R"%string))) (EVar "Rs"%string))]));([(PVar "_10"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "case_clause"%string));(EVar "_10"%string)])]))]));([(PVar "_11"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "case_clause"%string));(EVar "_11"%string)])]))]));([(PVar "_12"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "case_clause"%string));(EVar "_12"%string)])]))]));([(PVar "Y"%string);(PVar "X"%string);(PVar "Fun"%string);PNil;(PVar "R"%string);(PVar "Rs"%string);(PVar "S"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rufmergel"%string, 3)) [(ECons (ECons (EVar "S"%string) ENil) (ECons (ECons (EVar "Y"%string) (ECons (EVar "X"%string) (EVar "R"%string))) (EVar "Rs"%string)));ENil;(EVar "Fun"%string)]));([(PVar "_19"%string);(PVar "_18"%string);(PVar "_17"%string);(PVar "_16"%string);(PVar "_15"%string);(PVar "_14"%string);(PVar "_13"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_19"%string);(EVar "_18"%string);(EVar "_17"%string);(EVar "_16"%string);(EVar "_15"%string);(EVar "_14"%string);(EVar "_13"%string)])]))]) |};
          {| identifier := ("ufsplit_2"%string, 4) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string)]) [([(PVar "Y"%string);(PCons (PVar "Z"%string) (PVar "L"%string));(PVar "Fun"%string);(PVar "R"%string)], (ELit (Atom "true"%string)), (ECase (EApp (EVar "Fun"%string) [(EVar "Y"%string);(EVar "Z"%string)]) [([(PLit (Atom "true"%string))], (ELit (Atom "true"%string)), (ECase (EApp (EVar "Fun"%string) [(EVar "Z"%string);(EVar "Y"%string)]) [([(PLit (Atom "true"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("ufsplit_2"%string, 4)) [(EVar "Y"%string);(EVar "L"%string);(EVar "Fun"%string);(EVar "R"%string)]));([(PLit (Atom "false"%string))], (ELit (Atom "true"%string)), (ELet ["_4"%string] (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "R"%string);ENil]) (EApp (EFunId ("ufsplit_1"%string, 6)) [(EVar "Z"%string);(EVar "Y"%string);(EVar "Fun"%string);(EVar "L"%string);ENil;(ECons (EVar "_4"%string) ENil)])));([(PVar "_5"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "case_clause"%string));(EVar "_5"%string)])]))]));([(PLit (Atom "false"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("ufsplit_2"%string, 4)) [(EVar "Z"%string);(EVar "L"%string);(EVar "Fun"%string);(ECons (EVar "Y"%string) (EVar "R"%string))]));([(PVar "_6"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "case_clause"%string));(EVar "_6"%string)])]))]));([(PVar "Y"%string);PNil;(PVar "_Fun"%string);(PVar "R"%string)], (ELit (Atom "true"%string)), (ECons (EVar "Y"%string) (EVar "R"%string)));([(PVar "_10"%string);(PVar "_9"%string);(PVar "_8"%string);(PVar "_7"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_10"%string);(EVar "_9"%string);(EVar "_8"%string);(EVar "_7"%string)])]))]) |};
          {| identifier := ("ufmergel"%string, 3) ; varl := ["_0"%string;"_1"%string;"_2"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string)]) [([(PCons (PCons (PVar "H1"%string) (PVar "T1"%string)) (PCons (PVar "T2"%string) (PVar "L"%string)));(PVar "Acc"%string);(PVar "Fun"%string)], (ELit (Atom "true"%string)), (ELet ["_3"%string] (EApp (EFunId ("ufmerge2_2"%string, 5)) [(EVar "H1"%string);(EVar "T1"%string);(EVar "Fun"%string);(EVar "T2"%string);ENil]) (EApp (EFunId ("ufmergel"%string, 3)) [(EVar "L"%string);(ECons (EVar "_3"%string) (EVar "Acc"%string));(EVar "Fun"%string)])));([(PCons (PVar "L"%string) PNil);PNil;(PVar "_Fun"%string)], (ELit (Atom "true"%string)), (EVar "L"%string));([(PCons (PVar "L"%string) PNil);(PVar "Acc"%string);(PVar "Fun"%string)], (ELit (Atom "true"%string)), (ELet ["_4"%string] (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "L"%string);ENil]) (EApp (EFunId ("rufmergel"%string, 3)) [(ECons (EVar "_4"%string) (EVar "Acc"%string));ENil;(EVar "Fun"%string)])));([PNil;(PVar "Acc"%string);(PVar "Fun"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("rufmergel"%string, 3)) [(EVar "Acc"%string);ENil;(EVar "Fun"%string)]));([(PVar "_7"%string);(PVar "_6"%string);(PVar "_5"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_7"%string);(EVar "_6"%string);(EVar "_5"%string)])]))]) |};
          {| identifier := ("rufmergel"%string, 3) ; varl := ["_0"%string;"_1"%string;"_2"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string)]) [([(PCons (PCons (PVar "H2"%string) (PVar "T2"%string)) (PCons (PVar "T1"%string) (PVar "L"%string)));(PVar "Acc"%string);(PVar "Fun"%string)], (ELit (Atom "true"%string)), (ELet ["_3"%string] (EApp (EFunId ("rufmerge2_1"%string, 5)) [(EVar "T1"%string);(EVar "H2"%string);(EVar "Fun"%string);(EVar "T2"%string);ENil]) (EApp (EFunId ("rufmergel"%string, 3)) [(EVar "L"%string);(ECons (EVar "_3"%string) (EVar "Acc"%string));(EVar "Fun"%string)])));([(PCons (PVar "L"%string) PNil);(PVar "Acc"%string);(PVar "Fun"%string)], (ELit (Atom "true"%string)), (ELet ["_4"%string] (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "L"%string);ENil]) (EApp (EFunId ("ufmergel"%string, 3)) [(ECons (EVar "_4"%string) (EVar "Acc"%string));ENil;(EVar "Fun"%string)])));([PNil;(PVar "Acc"%string);(PVar "Fun"%string)], (ELit (Atom "true"%string)), (EApp (EFunId ("ufmergel"%string, 3)) [(EVar "Acc"%string);ENil;(EVar "Fun"%string)]));([(PVar "_7"%string);(PVar "_6"%string);(PVar "_5"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_7"%string);(EVar "_6"%string);(EVar "_5"%string)])]))]) |};
          {| identifier := ("ufmerge2_1"%string, 6) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string)]) [([(PCons (PVar "H1"%string) (PVar "T1"%string));(PVar "H2"%string);(PVar "Fun"%string);(PVar "T2"%string);(PVar "M"%string);(PVar "HdM"%string)], (ELit (Atom "true"%string)), (ECase (EApp (EVar "Fun"%string) [(EVar "H1"%string);(EVar "H2"%string)]) [([(PLit (Atom "true"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("ufmerge2_1"%string, 6)) [(EVar "T1"%string);(EVar "H2"%string);(EVar "Fun"%string);(EVar "T2"%string);(ECons (EVar "H1"%string) (EVar "M"%string));(EVar "H1"%string)]));([(PLit (Atom "false"%string))], (ELit (Atom "true"%string)), (ECase (EApp (EVar "Fun"%string) [(EVar "H2"%string);(EVar "HdM"%string)]) [([(PLit (Atom "true"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("ufmerge2_2"%string, 5)) [(EVar "H1"%string);(EVar "T1"%string);(EVar "Fun"%string);(EVar "T2"%string);(EVar "M"%string)]));([(PLit (Atom "false"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("ufmerge2_2"%string, 5)) [(EVar "H1"%string);(EVar "T1"%string);(EVar "Fun"%string);(EVar "T2"%string);(ECons (EVar "H2"%string) (EVar "M"%string))]));([(PVar "_6"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "case_clause"%string));(EVar "_6"%string)])]))]));([(PVar "_7"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "case_clause"%string));(EVar "_7"%string)])]))]));([PNil;(PVar "H2"%string);(PVar "Fun"%string);(PVar "T2"%string);(PVar "M"%string);(PVar "HdM"%string)], (ELit (Atom "true"%string)), (ECase (EApp (EVar "Fun"%string) [(EVar "H2"%string);(EVar "HdM"%string)]) [([(PLit (Atom "true"%string))], (ELit (Atom "true"%string)), (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "T2"%string);(EVar "M"%string)]));([(PLit (Atom "false"%string))], (ELit (Atom "true"%string)), (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "T2"%string);(ECons (EVar "H2"%string) (EVar "M"%string))]));([(PVar "_8"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "case_clause"%string));(EVar "_8"%string)])]))]));([(PVar "_14"%string);(PVar "_13"%string);(PVar "_12"%string);(PVar "_11"%string);(PVar "_10"%string);(PVar "_9"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_14"%string);(EVar "_13"%string);(EVar "_12"%string);(EVar "_11"%string);(EVar "_10"%string);(EVar "_9"%string)])]))]) |};
          {| identifier := ("ufmerge2_2"%string, 5) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string)]) [([(PVar "H1"%string);(PVar "T1"%string);(PVar "Fun"%string);(PCons (PVar "H2"%string) (PVar "T2"%string));(PVar "M"%string)], (ELit (Atom "true"%string)), (ECase (EApp (EVar "Fun"%string) [(EVar "H1"%string);(EVar "H2"%string)]) [([(PLit (Atom "true"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("ufmerge2_1"%string, 6)) [(EVar "T1"%string);(EVar "H2"%string);(EVar "Fun"%string);(EVar "T2"%string);(ECons (EVar "H1"%string) (EVar "M"%string));(EVar "H1"%string)]));([(PLit (Atom "false"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("ufmerge2_2"%string, 5)) [(EVar "H1"%string);(EVar "T1"%string);(EVar "Fun"%string);(EVar "T2"%string);(ECons (EVar "H2"%string) (EVar "M"%string))]));([(PVar "_5"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "case_clause"%string));(EVar "_5"%string)])]))]));([(PVar "H1"%string);(PVar "T1"%string);(PVar "_Fun"%string);PNil;(PVar "M"%string)], (ELit (Atom "true"%string)), (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "T1"%string);(ECons (EVar "H1"%string) (EVar "M"%string))]));([(PVar "_10"%string);(PVar "_9"%string);(PVar "_8"%string);(PVar "_7"%string);(PVar "_6"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_10"%string);(EVar "_9"%string);(EVar "_8"%string);(EVar "_7"%string);(EVar "_6"%string)])]))]) |};
          {| identifier := ("rufmerge2_1"%string, 5) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string)]) [([(PCons (PVar "H1"%string) (PVar "T1"%string));(PVar "H2"%string);(PVar "Fun"%string);(PVar "T2"%string);(PVar "M"%string)], (ELit (Atom "true"%string)), (ECase (EApp (EVar "Fun"%string) [(EVar "H1"%string);(EVar "H2"%string)]) [([(PLit (Atom "true"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("rufmerge2_2"%string, 6)) [(EVar "H1"%string);(EVar "T1"%string);(EVar "Fun"%string);(EVar "T2"%string);(EVar "M"%string);(EVar "H2"%string)]));([(PLit (Atom "false"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("rufmerge2_1"%string, 5)) [(EVar "T1"%string);(EVar "H2"%string);(EVar "Fun"%string);(EVar "T2"%string);(ECons (EVar "H1"%string) (EVar "M"%string))]));([(PVar "_5"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "case_clause"%string));(EVar "_5"%string)])]))]));([PNil;(PVar "H2"%string);(PVar "_Fun"%string);(PVar "T2"%string);(PVar "M"%string)], (ELit (Atom "true"%string)), (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "T2"%string);(ECons (EVar "H2"%string) (EVar "M"%string))]));([(PVar "_10"%string);(PVar "_9"%string);(PVar "_8"%string);(PVar "_7"%string);(PVar "_6"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_10"%string);(EVar "_9"%string);(EVar "_8"%string);(EVar "_7"%string);(EVar "_6"%string)])]))]) |};
          {| identifier := ("rufmerge2_2"%string, 6) ; varl := ["_0"%string;"_1"%string;"_2"%string;"_3"%string;"_4"%string;"_5"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string);(EVar "_3"%string);(EVar "_4"%string);(EVar "_5"%string)]) [([(PVar "H1"%string);(PVar "T1"%string);(PVar "Fun"%string);(PCons (PVar "H2"%string) (PVar "T2"%string));(PVar "M"%string);(PVar "H2M"%string)], (ELit (Atom "true"%string)), (ECase (EApp (EVar "Fun"%string) [(EVar "H1"%string);(EVar "H2"%string)]) [([(PLit (Atom "true"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("rufmerge2_2"%string, 6)) [(EVar "H1"%string);(EVar "T1"%string);(EVar "Fun"%string);(EVar "T2"%string);(ECons (EVar "H2M"%string) (EVar "M"%string));(EVar "H2"%string)]));([(PLit (Atom "false"%string))], (ELit (Atom "true"%string)), (ECase (EApp (EVar "Fun"%string) [(EVar "H2M"%string);(EVar "H1"%string)]) [([(PLit (Atom "true"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("rufmerge2_1"%string, 5)) [(EVar "T1"%string);(EVar "H2"%string);(EVar "Fun"%string);(EVar "T2"%string);(ECons (EVar "H1"%string) (EVar "M"%string))]));([(PLit (Atom "false"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("rufmerge2_1"%string, 5)) [(EVar "T1"%string);(EVar "H2"%string);(EVar "Fun"%string);(EVar "T2"%string);(ECons (EVar "H1"%string) (ECons (EVar "H2M"%string) (EVar "M"%string)))]));([(PVar "_6"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "case_clause"%string));(EVar "_6"%string)])]))]));([(PVar "_7"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "case_clause"%string));(EVar "_7"%string)])]))]));([(PVar "H1"%string);(PVar "T1"%string);(PVar "Fun"%string);PNil;(PVar "M"%string);(PVar "H2M"%string)], (ELit (Atom "true"%string)), (ECase (EApp (EVar "Fun"%string) [(EVar "H2M"%string);(EVar "H1"%string)]) [([(PLit (Atom "true"%string))], (ELit (Atom "true"%string)), (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "T1"%string);(ECons (EVar "H1"%string) (EVar "M"%string))]));([(PLit (Atom "false"%string))], (ELit (Atom "true"%string)), (ECall (ELit (Atom "lists"%string)) (ELit (Atom "reverse"%string)) [(EVar "T1"%string);(ECons (EVar "H1"%string) (ECons (EVar "H2M"%string) (EVar "M"%string)))]));([(PVar "_8"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "case_clause"%string));(EVar "_8"%string)])]))]));([(PVar "_14"%string);(PVar "_13"%string);(PVar "_12"%string);(PVar "_11"%string);(PVar "_10"%string);(PVar "_9"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_14"%string);(EVar "_13"%string);(EVar "_12"%string);(EVar "_11"%string);(EVar "_10"%string);(EVar "_9"%string)])]))]) |};
          {| identifier := ("uniq"%string, 1) ; varl := ["_0"%string]; body := (EApp (EFunId ("uniq_1"%string, 2)) [(EVar "_0"%string);(EMap [])]) |};
          {| identifier := ("uniq_1"%string, 2) ; varl := ["_0"%string;"_1"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string)]) [([(PCons (PVar "X"%string) (PVar "Xs"%string));(PVar "M"%string)], (ELit (Atom "true"%string)), (ECase (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_map_key"%string)) [(EVar "X"%string);(EVar "M"%string)]) [([(PLit (Atom "true"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("uniq_1"%string, 2)) [(EVar "Xs"%string);(EVar "M"%string)]));([(PLit (Atom "false"%string))], (ELit (Atom "true"%string)), (ECase (EValues []) [([], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_map"%string)) [(EVar "M"%string)]), (ELet ["_2"%string] (EMap [((EVar "X"%string), (ELit (Atom "true"%string)))]) (ELet ["_3"%string] (EApp (EFunId ("uniq_1"%string, 2)) [(EVar "Xs"%string);(EVar "_2"%string)]) (ECons (EVar "X"%string) (EVar "_3"%string)))));([], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "badmap"%string));(EVar "M"%string)])]))]));([(PVar "_4"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "case_clause"%string));(EVar "_4"%string)])]))]));([PNil;(PVar "_7"%string)], (ELit (Atom "true"%string)), ENil);([(PVar "_6"%string);(PVar "_5"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_6"%string);(EVar "_5"%string)])]))]) |};
          {| identifier := ("uniq"%string, 2) ; varl := ["_0"%string;"_1"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string)]) [([(PVar "F"%string);(PVar "L"%string)], (ETry (ELet ["_2"%string] (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_function"%string)) [(EVar "F"%string);(ELit (Integer (1)))]) (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "=:="%string)) [(EVar "_2"%string);(ELit (Atom "true"%string))])) ["Try"%string] (EVar "Try"%string) ["T"%string;"R"%string] (ELit (Atom "false"%string))), (EApp (EFunId ("uniq_2"%string, 3)) [(EVar "L"%string);(EVar "F"%string);(EMap [])]));([(PVar "_4"%string);(PVar "_3"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_4"%string);(EVar "_3"%string)])]))]) |};
          {| identifier := ("uniq_2"%string, 3) ; varl := ["_0"%string;"_1"%string;"_2"%string]; body := (ECase (EValues [(EVar "_0"%string);(EVar "_1"%string);(EVar "_2"%string)]) [([(PCons (PVar "X"%string) (PVar "Xs"%string));(PVar "F"%string);(PVar "M"%string)], (ELit (Atom "true"%string)), (ELet ["Key"%string] (EApp (EVar "F"%string) [(EVar "X"%string)]) (ECase (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_map_key"%string)) [(EVar "Key"%string);(EVar "M"%string)]) [([(PLit (Atom "true"%string))], (ELit (Atom "true"%string)), (EApp (EFunId ("uniq_2"%string, 3)) [(EVar "Xs"%string);(EVar "F"%string);(EVar "M"%string)]));([(PLit (Atom "false"%string))], (ELit (Atom "true"%string)), (ECase (EValues []) [([], (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "is_map"%string)) [(EVar "M"%string)]), (ELet ["_4"%string] (EMap [((EVar "Key"%string), (ELit (Atom "true"%string)))]) (ELet ["_5"%string] (EApp (EFunId ("uniq_2"%string, 3)) [(EVar "Xs"%string);(EVar "F"%string);(EVar "_4"%string)]) (ECons (EVar "X"%string) (EVar "_5"%string)))));([], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "badmap"%string));(EVar "M"%string)])]))]));([(PVar "_6"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "case_clause"%string));(EVar "_6"%string)])]))])));([PNil;(PVar "_10"%string);(PVar "_11"%string)], (ELit (Atom "true"%string)), ENil);([(PVar "_9"%string);(PVar "_8"%string);(PVar "_7"%string)], (ELit (Atom "true"%string)), (EPrimOp "match_fail"%string [(ETuple [(ELit (Atom "function_clause"%string));(EVar "_9"%string);(EVar "_8"%string);(EVar "_7"%string)])]))]) |};
          {| identifier := ("module_info"%string, 0) ; varl := []; body := (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "get_module_info"%string)) [(ELit (Atom "lists"%string))]) |};
          {| identifier := ("module_info"%string, 1) ; varl := ["_0"%string]; body := (ECall (ELit (Atom "erlang"%string)) (ELit (Atom "get_module_info"%string)) [(ELit (Atom "lists"%string));(EVar "_0"%string)]) |}
      ] 
    |}
  ] 
.


Definition valid_modules (ml : list ErlModule) : Prop := get_module "erlang"%string ml = None /\ get_module "io"%string ml = None /\ get_module "lists"%string ml = None.
Definition empty_modules (ml : list ErlModule) : Prop := ml = [].

 

Lemma module_concat1: 
  forall mname modules1 modules2, 
    get_module mname (modules1) = None ->
    get_module mname (modules2) = None -> 
    get_module mname (modules1 ++ modules2) = None .
Proof.
intros.
induction modules1.
  - simpl. exact H0.
  - inversion H. simpl. destruct ((name a =? mname)%string) eqn: A.
    -- auto.
    --  rewrite H2. apply (IHmodules1) in H2. rewrite H2. auto.
  
Qed.

Lemma module_concat2: 
  forall mname modules1 modules2, 
    get_module mname (modules1 ++ modules2) = None 
    ->
    get_module mname (modules1) = None /\
    get_module mname (modules2) = None
    .
Proof.
intros.
induction modules1.
  - auto.
  - simpl. inversion H. destruct ((name a =? mname)%string) eqn: A.
    -- congruence.
    -- rewrite H1. apply IHmodules1 in H1. auto. 
Qed.

Lemma module_rhs :
  forall mname modules1 modules2,
    get_module mname (modules2) = None ->
    get_module mname (modules1 ++ modules2) = get_module mname (modules1).
Proof.
  intros.
  induction modules1.
  - auto.
  - simpl. destruct ((name a =? mname)%string) eqn: A.
    -- auto.
    -- rewrite IHmodules1. auto.
Qed.

Lemma module_lhs :
  forall mname modules1 modules2,
    get_module mname (modules1) = None ->
    get_module mname (modules1 ++ modules2) = get_module mname (modules2).
Proof.
  intros.
  induction modules1.
  - auto.
  - inversion H. simpl. destruct ((name a =? mname)%string) eqn: A.
    -- congruence.
    -- auto. 
Qed.
